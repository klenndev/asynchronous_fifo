`ifndef CLK_CYCLE_SND
`define CLK_CYCLE_SND 5
`endif

`ifndef CLK_CYCLE_RCV
`define CLK_CYCLE_RCV 10
`endif


* cell custom_sram_1r1w_32_256_freepdk45
* pin addr0[0]
* pin addr0[1]
* pin din0[0]
* pin din0[1]
* pin din0[2]
* pin din0[3]
* pin din0[4]
* pin din0[5]
* pin din0[6]
* pin din0[7]
* pin din0[8]
* pin din0[9]
* pin din0[10]
* pin din0[11]
* pin din0[12]
* pin din0[13]
* pin din0[14]
* pin din0[15]
* pin din0[16]
* pin din0[17]
* pin din0[18]
* pin din0[19]
* pin din0[20]
* pin din0[21]
* pin din0[22]
* pin din0[23]
* pin din0[24]
* pin din0[25]
* pin din0[26]
* pin din0[27]
* pin din0[28]
* pin din0[29]
* pin din0[30]
* pin din0[31]
* pin csb0
* pin clk0
* pin addr1[7]
* pin addr1[6]
* pin addr1[5]
* pin addr1[4]
* pin addr1[3]
* pin addr1[2]
* pin addr0[5]
* pin addr0[4]
* pin addr0[3]
* pin addr0[2]
* pin addr0[6]
* pin addr0[7]
* pin dout1[0]
* pin dout1[1]
* pin dout1[2]
* pin dout1[3]
* pin dout1[4]
* pin dout1[5]
* pin dout1[6]
* pin dout1[7]
* pin dout1[8]
* pin dout1[9]
* pin dout1[10]
* pin dout1[11]
* pin dout1[12]
* pin dout1[13]
* pin dout1[14]
* pin dout1[15]
* pin dout1[16]
* pin dout1[17]
* pin dout1[18]
* pin dout1[19]
* pin dout1[20]
* pin dout1[21]
* pin dout1[22]
* pin dout1[23]
* pin dout1[24]
* pin dout1[25]
* pin dout1[26]
* pin dout1[27]
* pin dout1[28]
* pin dout1[29]
* pin dout1[30]
* pin dout1[31]
* pin clk1
* pin csb1
* pin addr1[1]
* pin addr1[0]
* pin NWELL
* pin BULK,PWELL
.SUBCKT custom_sram_1r1w_32_256_freepdk45 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 39 40 42 46 49
+ 52 55 56 57 58 63 65 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89
+ 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108
* net 2 addr0[0]
* net 3 addr0[1]
* net 4 din0[0]
* net 5 din0[1]
* net 6 din0[2]
* net 7 din0[3]
* net 8 din0[4]
* net 9 din0[5]
* net 10 din0[6]
* net 11 din0[7]
* net 12 din0[8]
* net 13 din0[9]
* net 14 din0[10]
* net 15 din0[11]
* net 16 din0[12]
* net 17 din0[13]
* net 18 din0[14]
* net 19 din0[15]
* net 20 din0[16]
* net 21 din0[17]
* net 22 din0[18]
* net 23 din0[19]
* net 24 din0[20]
* net 25 din0[21]
* net 26 din0[22]
* net 27 din0[23]
* net 28 din0[24]
* net 29 din0[25]
* net 30 din0[26]
* net 31 din0[27]
* net 32 din0[28]
* net 33 din0[29]
* net 34 din0[30]
* net 35 din0[31]
* net 36 csb0
* net 37 clk0
* net 39 addr1[7]
* net 40 addr1[6]
* net 42 addr1[5]
* net 46 addr1[4]
* net 49 addr1[3]
* net 52 addr1[2]
* net 55 addr0[5]
* net 56 addr0[4]
* net 57 addr0[3]
* net 58 addr0[2]
* net 63 addr0[6]
* net 65 addr0[7]
* net 71 dout1[0]
* net 72 dout1[1]
* net 73 dout1[2]
* net 74 dout1[3]
* net 75 dout1[4]
* net 76 dout1[5]
* net 77 dout1[6]
* net 78 dout1[7]
* net 79 dout1[8]
* net 80 dout1[9]
* net 81 dout1[10]
* net 82 dout1[11]
* net 83 dout1[12]
* net 84 dout1[13]
* net 85 dout1[14]
* net 86 dout1[15]
* net 87 dout1[16]
* net 88 dout1[17]
* net 89 dout1[18]
* net 90 dout1[19]
* net 91 dout1[20]
* net 92 dout1[21]
* net 93 dout1[22]
* net 94 dout1[23]
* net 95 dout1[24]
* net 96 dout1[25]
* net 97 dout1[26]
* net 98 dout1[27]
* net 99 dout1[28]
* net 100 dout1[29]
* net 101 dout1[30]
* net 102 dout1[31]
* net 103 clk1
* net 104 csb1
* net 105 addr1[1]
* net 106 addr1[0]
* net 107 NWELL
* net 108 BULK,PWELL
* cell instance $1 r0 *1 0.07,4.025
X$1 1 36 50 38 45 43 37 107 108
+ custom_sram_1r1w_32_256_freepdk45_control_logic_w
* cell instance $2 r0 *1 15.83,48.615
X$2 58 59 57 60 56 61 55 62 63 64 65 67 1 107 108
+ custom_sram_1r1w_32_256_freepdk45_row_addr_dff
* cell instance $3 r0 *1 27.27,0
X$3 1 4 133 5 142 6 139 7 113 8 136 9 132 10 125 11 141 12 138 13 115 14 130 15
+ 135 16 128 17 131 18 126 19 124 20 140 21 123 22 122 23 121 24 120 25 119 26
+ 118 27 117 28 137 29 116 30 114 31 129 32 112 33 134 34 127 35 111 107 108
+ custom_sram_1r1w_32_256_freepdk45_data_dff
* cell instance $4 r0 *1 21.55,0
X$4 2 144 3 143 1 107 108 custom_sram_1r1w_32_256_freepdk45_col_addr_dff
* cell instance $44 r0 *1 18.97,8.35
X$44 144 133 142 139 113 136 132 125 141 138 115 130 135 128 131 126 124 140
+ 123 122 121 120 119 118 117 137 116 114 129 112 134 127 111 38 143 43 45 59
+ 60 61 62 64 67 50 66 41 44 48 47 51 54 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 68 69 110 109
+ 107 108 custom_sram_1r1w_32_256_freepdk45_bank
* cell instance $47 r180 *1 269.275,24.695
X$47 52 54 49 51 46 47 42 48 40 44 39 41 53 107 108
+ custom_sram_1r1w_32_256_freepdk45_row_addr_dff
* cell instance $70 r180 *1 285.035,138.395
X$70 53 104 66 68 70 69 103 107 108
+ custom_sram_1r1w_32_256_freepdk45_control_logic_r
* cell instance $71 r180 *1 260.695,139.77
X$71 106 109 105 110 53 107 108 custom_sram_1r1w_32_256_freepdk45_col_addr_dff
.ENDS custom_sram_1r1w_32_256_freepdk45

* cell custom_sram_1r1w_32_256_freepdk45_row_addr_dff
* pin din_0
* pin dout_0
* pin din_1
* pin dout_1
* pin din_2
* pin dout_2
* pin din_3
* pin dout_3
* pin din_4
* pin dout_4
* pin din_5
* pin dout_5
* pin clk
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_row_addr_dff 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15
* net 1 din_0
* net 2 dout_0
* net 3 din_1
* net 4 dout_1
* net 5 din_2
* net 6 dout_2
* net 7 din_3
* net 8 dout_3
* net 9 din_4
* net 10 dout_4
* net 11 din_5
* net 12 dout_5
* net 13 clk
* net 14 vdd
* net 15 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 13 14 15 dff
* cell instance $2 m0 *1 0,4.94
X$2 4 3 13 14 15 dff
* cell instance $3 r0 *1 0,4.94
X$3 6 5 13 14 15 dff
* cell instance $4 m0 *1 0,9.88
X$4 8 7 13 14 15 dff
* cell instance $5 r0 *1 0,9.88
X$5 10 9 13 14 15 dff
* cell instance $6 m0 *1 0,14.82
X$6 12 11 13 14 15 dff
.ENDS custom_sram_1r1w_32_256_freepdk45_row_addr_dff

* cell custom_sram_1r1w_32_256_freepdk45_data_dff
* pin clk
* pin din_0
* pin dout_0
* pin din_1
* pin dout_1
* pin din_2
* pin dout_2
* pin din_3
* pin dout_3
* pin din_4
* pin dout_4
* pin din_5
* pin dout_5
* pin din_6
* pin dout_6
* pin din_7
* pin dout_7
* pin din_8
* pin dout_8
* pin din_9
* pin dout_9
* pin din_10
* pin dout_10
* pin din_11
* pin dout_11
* pin din_12
* pin dout_12
* pin din_13
* pin dout_13
* pin din_14
* pin dout_14
* pin din_15
* pin dout_15
* pin din_16
* pin dout_16
* pin din_17
* pin dout_17
* pin din_18
* pin dout_18
* pin din_19
* pin dout_19
* pin din_20
* pin dout_20
* pin din_21
* pin dout_21
* pin din_22
* pin dout_22
* pin din_23
* pin dout_23
* pin din_24
* pin dout_24
* pin din_25
* pin dout_25
* pin din_26
* pin dout_26
* pin din_27
* pin dout_27
* pin din_28
* pin dout_28
* pin din_29
* pin dout_29
* pin din_30
* pin dout_30
* pin din_31
* pin dout_31
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_data_dff 1 2 3 4 5 6 7 8 9 10 11 12
+ 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38
+ 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64
+ 65 66 67
* net 1 clk
* net 2 din_0
* net 3 dout_0
* net 4 din_1
* net 5 dout_1
* net 6 din_2
* net 7 dout_2
* net 8 din_3
* net 9 dout_3
* net 10 din_4
* net 11 dout_4
* net 12 din_5
* net 13 dout_5
* net 14 din_6
* net 15 dout_6
* net 16 din_7
* net 17 dout_7
* net 18 din_8
* net 19 dout_8
* net 20 din_9
* net 21 dout_9
* net 22 din_10
* net 23 dout_10
* net 24 din_11
* net 25 dout_11
* net 26 din_12
* net 27 dout_12
* net 28 din_13
* net 29 dout_13
* net 30 din_14
* net 31 dout_14
* net 32 din_15
* net 33 dout_15
* net 34 din_16
* net 35 dout_16
* net 36 din_17
* net 37 dout_17
* net 38 din_18
* net 39 dout_18
* net 40 din_19
* net 41 dout_19
* net 42 din_20
* net 43 dout_20
* net 44 din_21
* net 45 dout_21
* net 46 din_22
* net 47 dout_22
* net 48 din_23
* net 49 dout_23
* net 50 din_24
* net 51 dout_24
* net 52 din_25
* net 53 dout_25
* net 54 din_26
* net 55 dout_26
* net 56 din_27
* net 57 dout_27
* net 58 din_28
* net 59 dout_28
* net 60 din_29
* net 61 dout_29
* net 62 din_30
* net 63 dout_30
* net 64 din_31
* net 65 dout_31
* net 66 vdd
* net 67 gnd
* cell instance $1 r0 *1 88.66,0
X$1 65 64 1 66 67 dff
* cell instance $2 r0 *1 85.8,0
X$2 63 62 1 66 67 dff
* cell instance $3 r0 *1 82.94,0
X$3 61 60 1 66 67 dff
* cell instance $4 r0 *1 80.08,0
X$4 59 58 1 66 67 dff
* cell instance $5 r0 *1 77.22,0
X$5 57 56 1 66 67 dff
* cell instance $6 r0 *1 74.36,0
X$6 55 54 1 66 67 dff
* cell instance $7 r0 *1 71.5,0
X$7 53 52 1 66 67 dff
* cell instance $8 r0 *1 68.64,0
X$8 51 50 1 66 67 dff
* cell instance $9 r0 *1 65.78,0
X$9 49 48 1 66 67 dff
* cell instance $10 r0 *1 62.92,0
X$10 47 46 1 66 67 dff
* cell instance $11 r0 *1 60.06,0
X$11 45 44 1 66 67 dff
* cell instance $12 r0 *1 57.2,0
X$12 43 42 1 66 67 dff
* cell instance $13 r0 *1 54.34,0
X$13 41 40 1 66 67 dff
* cell instance $14 r0 *1 51.48,0
X$14 39 38 1 66 67 dff
* cell instance $15 r0 *1 48.62,0
X$15 37 36 1 66 67 dff
* cell instance $16 r0 *1 45.76,0
X$16 35 34 1 66 67 dff
* cell instance $17 r0 *1 2.86,0
X$17 5 4 1 66 67 dff
* cell instance $18 r0 *1 5.72,0
X$18 7 6 1 66 67 dff
* cell instance $19 r0 *1 8.58,0
X$19 9 8 1 66 67 dff
* cell instance $20 r0 *1 11.44,0
X$20 11 10 1 66 67 dff
* cell instance $21 r0 *1 14.3,0
X$21 13 12 1 66 67 dff
* cell instance $22 r0 *1 17.16,0
X$22 15 14 1 66 67 dff
* cell instance $23 r0 *1 20.02,0
X$23 17 16 1 66 67 dff
* cell instance $24 r0 *1 22.88,0
X$24 19 18 1 66 67 dff
* cell instance $25 r0 *1 25.74,0
X$25 21 20 1 66 67 dff
* cell instance $26 r0 *1 28.6,0
X$26 23 22 1 66 67 dff
* cell instance $27 r0 *1 31.46,0
X$27 25 24 1 66 67 dff
* cell instance $28 r0 *1 34.32,0
X$28 27 26 1 66 67 dff
* cell instance $29 r0 *1 37.18,0
X$29 29 28 1 66 67 dff
* cell instance $30 r0 *1 40.04,0
X$30 31 30 1 66 67 dff
* cell instance $31 r0 *1 0,0
X$31 3 2 1 66 67 dff
* cell instance $32 r0 *1 42.9,0
X$32 33 32 1 66 67 dff
.ENDS custom_sram_1r1w_32_256_freepdk45_data_dff

* cell custom_sram_1r1w_32_256_freepdk45_control_logic_w
* pin clk_buf
* pin csb
* pin wl_en
* pin w_en
* pin rbl_bl
* pin p_en_bar
* pin clk
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_control_logic_w 7 9 10 11 12 13 14 15
+ 16
* net 7 clk_buf
* net 9 csb
* net 10 wl_en
* net 11 w_en
* net 12 rbl_bl
* net 13 p_en_bar
* net 14 clk
* net 15 vdd
* net 16 gnd
* cell instance $1 r0 *1 6.105,9.88
X$1 6 4 1 15 16 custom_sram_1r1w_32_256_freepdk45_pnand2_1
* cell instance $2 r0 *1 7.0075,9.88
X$2 13 1 15 16 custom_sram_1r1w_32_256_freepdk45_pdriver_5
* cell instance $3 m0 *1 6.7925,4.94
X$3 5 2 8 15 16 custom_sram_1r1w_32_256_freepdk45_pand2_0
* cell instance $4 m0 *1 6.105,4.94
X$4 7 2 15 16 custom_sram_1r1w_32_256_freepdk45_pinv_4
* cell instance $5 m0 *1 6.105,9.88
X$5 11 8 3 5 15 16 custom_sram_1r1w_32_256_freepdk45_pand3
* cell instance $8 m0 *1 6.105,14.82
X$8 4 3 15 16 custom_sram_1r1w_32_256_freepdk45_pinv_4
* cell instance $11 m0 *1 0,32.11
X$11 4 12 15 16 custom_sram_1r1w_32_256_freepdk45_delay_chain
* cell instance $16 r0 *1 6.105,14.82
X$16 10 5 15 16 custom_sram_1r1w_32_256_freepdk45_pdriver_2
* cell instance $23 r0 *1 6.105,4.94
X$23 6 7 8 15 16 custom_sram_1r1w_32_256_freepdk45_pand2_0
* cell instance $28 r0 *1 0,0
X$28 9 8 7 15 16 custom_sram_1r1w_32_256_freepdk45_dff_buf_array
* cell instance $34 r0 *1 6.105,0
X$34 7 14 15 16 custom_sram_1r1w_32_256_freepdk45_pdriver_1
.ENDS custom_sram_1r1w_32_256_freepdk45_control_logic_w

* cell custom_sram_1r1w_32_256_freepdk45_control_logic_r
* pin clk_buf
* pin csb
* pin wl_en
* pin s_en
* pin rbl_bl
* pin p_en_bar
* pin clk
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_control_logic_r 6 8 9 10 11 12 13 14
+ 15
* net 6 clk_buf
* net 8 csb
* net 9 wl_en
* net 10 s_en
* net 11 rbl_bl
* net 12 p_en_bar
* net 13 clk
* net 14 vdd
* net 15 gnd
* cell instance $1 r0 *1 7.0075,9.88
X$1 12 1 14 15 custom_sram_1r1w_32_256_freepdk45_pdriver_5
* cell instance $2 r0 *1 6.105,9.88
X$2 5 3 1 14 15 custom_sram_1r1w_32_256_freepdk45_pnand2_1
* cell instance $3 m0 *1 6.7925,4.94
X$3 4 2 7 14 15 custom_sram_1r1w_32_256_freepdk45_pand2_0
* cell instance $4 m0 *1 6.105,4.94
X$4 6 2 14 15 custom_sram_1r1w_32_256_freepdk45_pinv_4
* cell instance $5 m0 *1 6.105,9.88
X$5 10 3 4 7 14 15 custom_sram_1r1w_32_256_freepdk45_pand3_0
* cell instance $6 m0 *1 0,32.11
X$6 3 11 14 15 custom_sram_1r1w_32_256_freepdk45_delay_chain
* cell instance $11 m0 *1 6.105,14.82
X$11 9 4 14 15 custom_sram_1r1w_32_256_freepdk45_pdriver_2
* cell instance $18 r0 *1 6.105,4.94
X$18 5 6 7 14 15 custom_sram_1r1w_32_256_freepdk45_pand2_0
* cell instance $22 r0 *1 0,0
X$22 8 7 6 14 15 custom_sram_1r1w_32_256_freepdk45_dff_buf_array
* cell instance $25 r0 *1 6.105,0
X$25 6 13 14 15 custom_sram_1r1w_32_256_freepdk45_pdriver_1
.ENDS custom_sram_1r1w_32_256_freepdk45_control_logic_r

* cell custom_sram_1r1w_32_256_freepdk45_col_addr_dff
* pin din_0
* pin dout_0
* pin din_1
* pin dout_1
* pin clk
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_col_addr_dff 1 2 3 4 5 6 7
* net 1 din_0
* net 2 dout_0
* net 3 din_1
* net 4 dout_1
* net 5 clk
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 5 6 7 dff
* cell instance $2 r0 *1 2.86,0
X$2 4 3 5 6 7 dff
.ENDS custom_sram_1r1w_32_256_freepdk45_col_addr_dff

* cell custom_sram_1r1w_32_256_freepdk45_bank
* pin addr0_0
* pin din0_0
* pin din0_1
* pin din0_2
* pin din0_3
* pin din0_4
* pin din0_5
* pin din0_6
* pin din0_7
* pin din0_8
* pin din0_9
* pin din0_10
* pin din0_11
* pin din0_12
* pin din0_13
* pin din0_14
* pin din0_15
* pin din0_16
* pin din0_17
* pin din0_18
* pin din0_19
* pin din0_20
* pin din0_21
* pin din0_22
* pin din0_23
* pin din0_24
* pin din0_25
* pin din0_26
* pin din0_27
* pin din0_28
* pin din0_29
* pin din0_30
* pin din0_31
* pin w_en0
* pin addr0_1
* pin p_en_bar0
* pin rbl_bl_0_0
* pin addr0_2
* pin addr0_3
* pin addr0_4
* pin addr0_5
* pin addr0_6
* pin addr0_7
* pin wl_en0
* pin wl_en1
* pin addr1_7
* pin addr1_6
* pin addr1_5
* pin addr1_4
* pin addr1_3
* pin addr1_2
* pin rbl_bl_1_1
* pin dout1_0
* pin dout1_1
* pin dout1_2
* pin dout1_3
* pin dout1_4
* pin dout1_5
* pin dout1_6
* pin dout1_7
* pin dout1_8
* pin dout1_9
* pin dout1_10
* pin dout1_11
* pin dout1_12
* pin dout1_13
* pin dout1_14
* pin dout1_15
* pin dout1_16
* pin dout1_17
* pin dout1_18
* pin dout1_19
* pin dout1_20
* pin dout1_21
* pin dout1_22
* pin dout1_23
* pin dout1_24
* pin dout1_25
* pin dout1_26
* pin dout1_27
* pin dout1_28
* pin dout1_29
* pin dout1_30
* pin dout1_31
* pin s_en1
* pin p_en_bar1
* pin addr1_1
* pin addr1_0
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_bank 1 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 39 41 299
+ 300 301 302 303 304 305 436 437 438 439 440 441 442 699 701 702 703 704 705
+ 706 707 708 709 710 711 712 713 714 715 716 717 718 719 720 721 722 723 724
+ 725 726 727 728 729 730 731 732 737 738 739 740 741 742
* net 1 addr0_0
* net 4 din0_0
* net 5 din0_1
* net 6 din0_2
* net 7 din0_3
* net 8 din0_4
* net 9 din0_5
* net 10 din0_6
* net 11 din0_7
* net 12 din0_8
* net 13 din0_9
* net 14 din0_10
* net 15 din0_11
* net 16 din0_12
* net 17 din0_13
* net 18 din0_14
* net 19 din0_15
* net 20 din0_16
* net 21 din0_17
* net 22 din0_18
* net 23 din0_19
* net 24 din0_20
* net 25 din0_21
* net 26 din0_22
* net 27 din0_23
* net 28 din0_24
* net 29 din0_25
* net 30 din0_26
* net 31 din0_27
* net 32 din0_28
* net 33 din0_29
* net 34 din0_30
* net 35 din0_31
* net 36 w_en0
* net 37 addr0_1
* net 39 p_en_bar0
* net 41 rbl_bl_0_0
* net 299 addr0_2
* net 300 addr0_3
* net 301 addr0_4
* net 302 addr0_5
* net 303 addr0_6
* net 304 addr0_7
* net 305 wl_en0
* net 436 wl_en1
* net 437 addr1_7
* net 438 addr1_6
* net 439 addr1_5
* net 440 addr1_4
* net 441 addr1_3
* net 442 addr1_2
* net 699 rbl_bl_1_1
* net 701 dout1_0
* net 702 dout1_1
* net 703 dout1_2
* net 704 dout1_3
* net 705 dout1_4
* net 706 dout1_5
* net 707 dout1_6
* net 708 dout1_7
* net 709 dout1_8
* net 710 dout1_9
* net 711 dout1_10
* net 712 dout1_11
* net 713 dout1_12
* net 714 dout1_13
* net 715 dout1_14
* net 716 dout1_15
* net 717 dout1_16
* net 718 dout1_17
* net 719 dout1_18
* net 720 dout1_19
* net 721 dout1_20
* net 722 dout1_21
* net 723 dout1_22
* net 724 dout1_23
* net 725 dout1_24
* net 726 dout1_25
* net 727 dout1_26
* net 728 dout1_27
* net 729 dout1_28
* net 730 dout1_29
* net 731 dout1_30
* net 732 dout1_31
* net 737 s_en1
* net 738 p_en_bar1
* net 739 addr1_1
* net 740 addr1_0
* net 741 vdd
* net 742 gnd
* cell instance $1 r0 *1 4.585,0.1375
X$1 2 3 38 40 1 37 741 742 custom_sram_1r1w_32_256_freepdk45_column_decoder
* cell instance $2 m0 *1 12.71,13.105
X$2 41 42 43 44 45 46 47 48 49 51 52 53 54 55 56 57 58 59 61 62 63 64 65 66 67
+ 68 69 70 71 72 73 74 75 77 79 81 83 84 85 86 87 88 89 90 91 93 95 97 98 99
+ 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118
+ 119 120 121 123 124 125 126 127 128 129 130 131 133 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159
+ 160 161 162 163 164 165 166 167 168 169 171 172 173 174 175 176 177 178 179
+ 181 182 183 184 185 186 187 189 190 191 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 251 253 254 255 256 257 258 259 260 261
+ 262 263 264 265 267 269 270 271 272 273 274 275 277 279 280 281 282 283 284
+ 285 286 287 288 289 290 291 292 293 294 295 296 297 298 50 60 76 78 80 82 92
+ 94 96 122 132 134 170 39 180 188 192 210 250 252 266 268 276 278 4 5 6 7 8 9
+ 10 11 12 13 14 15 16 17 18 19 36 3 40 38 2 20 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 741 742 custom_sram_1r1w_32_256_freepdk45_port_data
* cell instance $11 r0 *1 12.71,13.105
X$11 356 359 363 366 369 345 344 332 329 335 337 321 311 308 315 318 326 323
+ 342 341 339 338 346 348 343 340 347 350 353 362 352 351 349 41 42 43 443 444
+ 44 45 445 446 46 47 447 448 48 49 449 450 50 51 451 452 52 53 453 454 54 55
+ 455 456 56 57 457 458 58 59 459 460 60 61 461 462 62 63 463 464 64 65 465 466
+ 66 67 467 468 68 69 469 470 70 71 471 472 72 73 473 474 74 75 475 476 76 77
+ 477 478 78 79 479 480 80 81 481 482 82 83 483 484 84 85 485 486 86 87 487 488
+ 88 89 489 490 90 91 491 492 92 93 493 494 94 95 495 496 96 97 497 498 98 99
+ 499 500 100 101 501 502 102 103 503 504 104 105 505 506 106 382 374 386 408
+ 371 380 427 378 383 423 405 396 393 395 373 392 399 397 398 394 379 385 404
+ 377 424 400 407 406 412 403 372 402 107 507 508 108 109 509 510 110 111 511
+ 512 112 113 513 514 114 115 515 516 116 117 517 518 118 119 519 520 120 121
+ 521 522 122 123 523 524 124 125 525 526 126 127 527 528 128 129 529 530 130
+ 131 531 532 132 133 533 534 134 135 535 536 136 137 537 538 138 139 539 540
+ 140 141 541 542 142 143 543 544 144 145 545 546 146 147 547 548 148 149 549
+ 550 150 151 551 552 152 153 553 554 154 155 555 556 156 157 557 558 158 159
+ 559 560 160 161 561 562 162 163 563 564 164 165 565 566 166 167 567 568 168
+ 169 569 570 170 171 571 572 172 173 573 574 174 175 575 576 176 177 577 578
+ 178 179 579 580 180 181 581 582 182 183 583 584 184 185 585 586 186 187 587
+ 588 188 189 589 590 190 191 591 592 192 193 593 594 194 195 595 596 196 197
+ 597 598 198 199 599 600 200 201 601 602 202 203 603 604 204 205 605 606 206
+ 207 607 608 208 209 609 610 210 211 611 612 212 213 613 614 214 215 615 616
+ 216 217 617 618 218 219 619 620 220 221 621 622 222 223 623 624 224 225 625
+ 626 226 227 627 628 228 229 629 630 230 231 631 632 232 233 633 634 234 235
+ 635 636 236 237 637 638 238 239 639 640 240 241 641 642 242 243 643 644 244
+ 245 645 646 246 247 647 648 248 249 649 650 250 251 651 652 252 253 653 654
+ 254 255 655 656 256 257 657 658 258 259 659 660 260 261 661 662 262 263 663
+ 664 264 265 665 666 266 267 667 668 268 269 669 670 270 271 671 672 272 273
+ 673 674 274 275 675 676 276 277 677 678 278 279 679 680 280 281 681 682 282
+ 283 683 684 284 285 685 686 286 287 687 688 288 289 689 690 290 291 691 692
+ 292 293 693 694 294 295 695 696 296 297 697 698 298 699 700 310 365 312 364
+ 313 354 355 361 336 357 334 316 314 317 370 306 319 360 307 368 320 309 367
+ 358 322 324 325 327 328 330 333 331 422 421 419 401 420 429 428 426 425 417
+ 391 390 389 388 387 376 384 381 418 416 415 414 413 411 410 409 435 434 375
+ 433 432 431 430 741 742 custom_sram_1r1w_32_256_freepdk45_global_bitcell_array
* cell instance $13 r0 *1 0,16.345
X$13 305 323 326 329 332 335 337 311 308 299 300 301 302 303 304 315 318 321
+ 356 359 363 366 369 345 344 343 340 347 350 353 362 352 351 349 348 346 338
+ 339 341 342 370 368 367 365 364 361 360 358 357 355 354 320 319 317 316 314
+ 306 307 309 310 312 313 336 334 333 331 330 328 327 325 324 322 741 742
+ custom_sram_1r1w_32_256_freepdk45_port_address
* cell instance $144 m90 *1 246.97,16.345
X$144 394 400 404 385 378 380 383 424 442 441 440 439 438 437 412 373 372 371
+ 374 408 423 427 386 382 379 377 407 406 403 402 396 393 395 397 398 399 392
+ 405 381 384 376 387 388 389 390 391 417 425 426 428 429 430 431 432 433 375
+ 434 435 409 410 411 413 414 415 416 418 419 420 421 436 422 401 741 742
+ custom_sram_1r1w_32_256_freepdk45_port_address_0
* cell instance $275 r0 *1 12.71,115.085
X$275 443 444 445 446 447 449 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 471 472 473 474 475 477 478 479 480 481 482 483
+ 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 511 512 513 515 516 517 518 519 520 521 522 523
+ 524 525 526 527 528 529 531 532 533 535 536 537 538 539 540 541 542 543 544
+ 545 546 547 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564
+ 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583
+ 584 585 587 588 589 590 591 592 593 595 596 597 598 599 600 601 602 603 604
+ 605 607 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625
+ 626 627 628 629 630 631 633 634 635 636 637 638 639 640 641 642 643 644 645
+ 646 647 648 649 650 651 652 653 654 655 656 657 659 660 661 663 664 665 666
+ 667 668 669 670 671 672 673 674 675 676 677 678 679 680 681 682 683 684 685
+ 686 687 688 689 690 691 692 693 694 695 696 697 698 699 700 448 450 470 476
+ 510 514 530 534 548 738 586 594 606 608 632 658 662 701 702 703 704 705 706
+ 707 708 709 710 711 712 713 714 715 716 737 734 733 735 736 717 718 719 720
+ 721 722 723 724 725 726 727 728 729 730 731 732 741 742
+ custom_sram_1r1w_32_256_freepdk45_port_data_0
* cell instance $277 r180 *1 242.385,128.0525
X$277 735 736 733 734 740 739 741 742
+ custom_sram_1r1w_32_256_freepdk45_column_decoder
.ENDS custom_sram_1r1w_32_256_freepdk45_bank

* cell custom_sram_1r1w_32_256_freepdk45_pand3
* pin Z
* pin A
* pin B
* pin C
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pand3 2 3 4 5 6 7
* net 2 Z
* net 3 A
* net 4 B
* net 5 C
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 0,0
X$1 3 4 5 1 6 7 custom_sram_1r1w_32_256_freepdk45_pnand3_0
* cell instance $2 r0 *1 0.965,0
X$2 2 1 6 7 custom_sram_1r1w_32_256_freepdk45_pdriver_3
.ENDS custom_sram_1r1w_32_256_freepdk45_pand3

* cell custom_sram_1r1w_32_256_freepdk45_pdriver_5
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pdriver_5 5 6 8 9
* net 5 Z
* net 6 A
* net 8 vdd
* net 9 gnd
* cell instance $1 r0 *1 1.375,0
X$1 1 2 8 9 custom_sram_1r1w_32_256_freepdk45_pinv_18
* cell instance $2 r0 *1 0.6875,0
X$2 7 1 8 9 custom_sram_1r1w_32_256_freepdk45_pinv_3
* cell instance $3 r0 *1 2.0625,0
X$3 2 3 8 9 custom_sram_1r1w_32_256_freepdk45_pinv_19
* cell instance $4 r0 *1 3.025,0
X$4 3 4 8 9 custom_sram_1r1w_32_256_freepdk45_pinv_20
* cell instance $5 r0 *1 4.8125,0
X$5 4 5 8 9 custom_sram_1r1w_32_256_freepdk45_pinv_21
* cell instance $6 r0 *1 0,0
X$6 6 7 8 9 custom_sram_1r1w_32_256_freepdk45_pinv_3
.ENDS custom_sram_1r1w_32_256_freepdk45_pdriver_5

* cell custom_sram_1r1w_32_256_freepdk45_pnand2_1
* pin A
* pin B
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pnand2_1 1 2 3 4 5
* net 1 A
* net 2 B
* net 3 Z
* net 4 vdd
* net 5 gnd
* device instance $1 r0 *1 0.2325,2.21 PMOS_VTG
M$1 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,2.21 PMOS_VTG
M$2 3 2 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.2325,0.215 NMOS_VTG
M$3 5 1 6 5 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $4 r0 *1 0.4475,0.215 NMOS_VTG
M$4 6 2 3 5 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS custom_sram_1r1w_32_256_freepdk45_pnand2_1

* cell custom_sram_1r1w_32_256_freepdk45_delay_chain
* pin out
* pin in
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_delay_chain 1 10 11 12
* net 1 out
* net 10 in
* net 11 vdd
* net 12 gnd
* cell instance $2 r0 *1 0.6875,19.76
X$2 1 37 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $5 r0 *1 1.375,19.76
X$5 1 36 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $8 r0 *1 2.0625,19.76
X$8 1 35 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $11 r0 *1 2.75,19.76
X$11 1 34 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $14 r0 *1 0,19.76
X$14 9 1 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $17 r0 *1 1.375,0
X$17 2 29 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $20 r0 *1 0.6875,0
X$20 2 46 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $23 m0 *1 0,4.94
X$23 2 3 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $25 r0 *1 2.0625,0
X$25 2 45 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $28 r0 *1 2.75,0
X$28 2 47 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $31 r0 *1 0,0
X$31 10 2 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $34 m0 *1 2.0625,4.94
X$34 3 22 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $37 r0 *1 0,4.94
X$37 3 4 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $39 m0 *1 2.75,4.94
X$39 3 23 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $42 m0 *1 0.6875,4.94
X$42 3 16 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $47 m0 *1 1.375,4.94
X$47 3 13 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $50 r0 *1 1.375,4.94
X$50 4 31 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $55 r0 *1 2.75,4.94
X$55 4 33 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $58 r0 *1 2.0625,4.94
X$58 4 32 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $61 m0 *1 0,9.88
X$61 4 5 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $63 r0 *1 0.6875,4.94
X$63 4 30 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $66 m0 *1 2.0625,9.88
X$66 5 15 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $69 r0 *1 0,9.88
X$69 5 6 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $71 m0 *1 0.6875,9.88
X$71 5 27 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $74 m0 *1 2.75,9.88
X$74 5 21 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $79 m0 *1 1.375,9.88
X$79 5 14 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $82 m0 *1 0,14.82
X$82 6 7 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $84 r0 *1 2.0625,9.88
X$84 6 43 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $87 r0 *1 0.6875,9.88
X$87 6 48 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $92 r0 *1 1.375,9.88
X$92 6 44 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $95 r0 *1 2.75,9.88
X$95 6 42 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $100 m0 *1 2.75,14.82
X$100 7 24 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $103 m0 *1 2.0625,14.82
X$103 7 25 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $106 m0 *1 0.6875,14.82
X$106 7 28 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $109 m0 *1 1.375,14.82
X$109 7 26 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $112 r0 *1 0,14.82
X$112 7 8 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $114 r0 *1 1.375,14.82
X$114 8 40 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $117 r0 *1 0.6875,14.82
X$117 8 41 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $120 r0 *1 2.0625,14.82
X$120 8 39 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $123 r0 *1 2.75,14.82
X$123 8 38 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $128 m0 *1 0,19.76
X$128 8 9 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $130 m0 *1 1.375,19.76
X$130 9 19 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $133 m0 *1 0.6875,19.76
X$133 9 20 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $136 m0 *1 2.0625,19.76
X$136 9 18 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
* cell instance $139 m0 *1 2.75,19.76
X$139 9 17 11 12 custom_sram_1r1w_32_256_freepdk45_pinv_22
.ENDS custom_sram_1r1w_32_256_freepdk45_delay_chain

* cell custom_sram_1r1w_32_256_freepdk45_pand3_0
* pin Z
* pin A
* pin B
* pin C
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pand3_0 2 3 4 5 6 7
* net 2 Z
* net 3 A
* net 4 B
* net 5 C
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 0.965,0
X$1 2 1 6 7 custom_sram_1r1w_32_256_freepdk45_pdriver_4
* cell instance $2 r0 *1 0,0
X$2 3 4 5 1 6 7 custom_sram_1r1w_32_256_freepdk45_pnand3_0
.ENDS custom_sram_1r1w_32_256_freepdk45_pand3_0

* cell custom_sram_1r1w_32_256_freepdk45_pdriver_2
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pdriver_2 2 3 4 5
* net 2 Z
* net 3 A
* net 4 vdd
* net 5 gnd
* cell instance $1 r0 *1 0,0
X$1 3 1 4 5 custom_sram_1r1w_32_256_freepdk45_pinv_14
* cell instance $2 r0 *1 1.2375,0
X$2 1 2 4 5 custom_sram_1r1w_32_256_freepdk45_pinv_15
.ENDS custom_sram_1r1w_32_256_freepdk45_pdriver_2

* cell custom_sram_1r1w_32_256_freepdk45_pand2_0
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pand2_0 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0.75,0
X$1 2 1 5 6 custom_sram_1r1w_32_256_freepdk45_pdriver_0
* cell instance $2 r0 *1 0,0
X$2 3 4 1 5 6 custom_sram_1r1w_32_256_freepdk45_pnand2_0
.ENDS custom_sram_1r1w_32_256_freepdk45_pand2_0

* cell custom_sram_1r1w_32_256_freepdk45_pdriver_1
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pdriver_1 5 6 8 9
* net 5 Z
* net 6 A
* net 8 vdd
* net 9 gnd
* cell instance $1 r0 *1 1.375,0
X$1 1 2 8 9 custom_sram_1r1w_32_256_freepdk45_pinv_10
* cell instance $2 r0 *1 0.6875,0
X$2 7 1 8 9 custom_sram_1r1w_32_256_freepdk45_pinv_3
* cell instance $3 r0 *1 2.0625,0
X$3 2 3 8 9 custom_sram_1r1w_32_256_freepdk45_pinv_11
* cell instance $4 r0 *1 3.3,0
X$4 3 4 8 9 custom_sram_1r1w_32_256_freepdk45_pinv_12
* cell instance $5 r0 *1 5.9125,0
X$5 4 5 8 9 custom_sram_1r1w_32_256_freepdk45_pinv_13
* cell instance $6 r0 *1 0,0
X$6 6 7 8 9 custom_sram_1r1w_32_256_freepdk45_pinv_3
.ENDS custom_sram_1r1w_32_256_freepdk45_pdriver_1

* cell custom_sram_1r1w_32_256_freepdk45_dff_buf_array
* pin din_0
* pin dout_bar_0
* pin clk
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_dff_buf_array 1 3 4 5 6
* net 1 din_0
* net 2 dout_0
* net 3 dout_bar_0
* net 4 clk
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0,0
X$1 3 2 4 1 5 6 custom_sram_1r1w_32_256_freepdk45_dff_buf_0
.ENDS custom_sram_1r1w_32_256_freepdk45_dff_buf_array

* cell custom_sram_1r1w_32_256_freepdk45_column_decoder
* pin out_0
* pin out_1
* pin out_2
* pin out_3
* pin in_0
* pin in_1
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_column_decoder 1 2 3 4 5 6 7 8
* net 1 out_0
* net 2 out_1
* net 3 out_2
* net 4 out_3
* net 5 in_0
* net 6 in_1
* net 7 vdd
* net 8 gnd
* cell instance $1 r0 *1 0,0
X$1 5 6 1 2 3 4 7 8
+ custom_sram_1r1w_32_256_freepdk45_hierarchical_predecode2x4_0
.ENDS custom_sram_1r1w_32_256_freepdk45_column_decoder

* cell custom_sram_1r1w_32_256_freepdk45_port_address_0
* pin wl_0
* pin wl_1
* pin wl_2
* pin wl_3
* pin wl_4
* pin wl_5
* pin wl_6
* pin wl_7
* pin addr_0
* pin addr_1
* pin addr_2
* pin addr_3
* pin addr_4
* pin addr_5
* pin wl_8
* pin wl_9
* pin wl_10
* pin wl_11
* pin wl_12
* pin wl_13
* pin wl_14
* pin wl_15
* pin wl_16
* pin wl_17
* pin wl_18
* pin wl_19
* pin wl_20
* pin wl_21
* pin wl_22
* pin wl_23
* pin wl_24
* pin wl_25
* pin wl_26
* pin wl_27
* pin wl_28
* pin wl_29
* pin wl_30
* pin wl_31
* pin wl_32
* pin wl_33
* pin wl_34
* pin wl_35
* pin wl_36
* pin wl_37
* pin wl_38
* pin wl_39
* pin wl_40
* pin wl_41
* pin wl_42
* pin wl_43
* pin wl_44
* pin wl_45
* pin wl_46
* pin wl_47
* pin wl_48
* pin wl_49
* pin wl_50
* pin wl_51
* pin wl_52
* pin wl_53
* pin wl_54
* pin wl_55
* pin wl_56
* pin wl_57
* pin wl_58
* pin wl_59
* pin wl_60
* pin wl_61
* pin wl_62
* pin wl_en
* pin wl_63
* pin rbl_wl
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_port_address_0 3 5 7 8 11 13 15 16 17
+ 18 19 20 21 22 25 26 29 31 33 34 36 38 41 42 45 46 49 50 53 54 57 58 61 62 65
+ 66 69 70 73 74 77 78 81 82 85 86 89 90 93 94 97 98 101 102 105 106 109 110
+ 113 114 117 118 121 122 125 126 129 130 133 134 135 136 137 138
* net 3 wl_0
* net 5 wl_1
* net 7 wl_2
* net 8 wl_3
* net 11 wl_4
* net 13 wl_5
* net 15 wl_6
* net 16 wl_7
* net 17 addr_0
* net 18 addr_1
* net 19 addr_2
* net 20 addr_3
* net 21 addr_4
* net 22 addr_5
* net 25 wl_8
* net 26 wl_9
* net 29 wl_10
* net 31 wl_11
* net 33 wl_12
* net 34 wl_13
* net 36 wl_14
* net 38 wl_15
* net 41 wl_16
* net 42 wl_17
* net 45 wl_18
* net 46 wl_19
* net 49 wl_20
* net 50 wl_21
* net 53 wl_22
* net 54 wl_23
* net 57 wl_24
* net 58 wl_25
* net 61 wl_26
* net 62 wl_27
* net 65 wl_28
* net 66 wl_29
* net 69 wl_30
* net 70 wl_31
* net 73 wl_32
* net 74 wl_33
* net 77 wl_34
* net 78 wl_35
* net 81 wl_36
* net 82 wl_37
* net 85 wl_38
* net 86 wl_39
* net 89 wl_40
* net 90 wl_41
* net 93 wl_42
* net 94 wl_43
* net 97 wl_44
* net 98 wl_45
* net 101 wl_46
* net 102 wl_47
* net 105 wl_48
* net 106 wl_49
* net 109 wl_50
* net 110 wl_51
* net 113 wl_52
* net 114 wl_53
* net 117 wl_54
* net 118 wl_55
* net 121 wl_56
* net 122 wl_57
* net 125 wl_58
* net 126 wl_59
* net 129 wl_60
* net 130 wl_61
* net 133 wl_62
* net 134 wl_en
* net 135 wl_63
* net 136 rbl_wl
* net 137 vdd
* net 138 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 18 17 4 6 9 10 14 12 19 20 21 22 23 28 27 24 30 35 32 40 39 37 43 44 47
+ 48 51 52 55 56 59 60 63 64 67 68 72 71 76 75 80 79 84 83 88 87 92 91 96 95
+ 100 99 104 103 108 107 112 111 116 115 120 119 124 123 128 127 132 131 137
+ 138 custom_sram_1r1w_32_256_freepdk45_hierarchical_decoder
* cell instance $2 r0 *1 8.515,0
X$2 1 3 2 5 4 7 6 8 10 11 9 13 12 15 14 16 23 25 24 26 28 29 27 31 30 33 32 34
+ 35 36 37 38 39 41 40 42 43 45 44 46 47 49 48 50 51 53 52 54 55 57 56 58 59 61
+ 60 62 63 65 64 66 67 69 68 134 70 72 73 74 71 76 77 78 75 80 81 82 79 84 85
+ 86 83 88 89 90 87 92 93 94 91 96 97 98 95 100 101 102 99 104 105 106 103 108
+ 109 110 107 112 113 114 111 116 117 118 115 120 121 122 119 124 125 126 123
+ 128 129 130 127 132 133 135 131 137 138
+ custom_sram_1r1w_32_256_freepdk45_wordline_driver_array
* cell instance $4 r0 *1 9.075,95.68
X$4 134 136 137 138 custom_sram_1r1w_32_256_freepdk45_pinv_2
.ENDS custom_sram_1r1w_32_256_freepdk45_port_address_0

* cell custom_sram_1r1w_32_256_freepdk45_port_address
* pin wl_en
* pin rbl_wl
* pin wl_0
* pin wl_1
* pin wl_2
* pin wl_3
* pin wl_4
* pin wl_5
* pin wl_6
* pin addr_0
* pin addr_1
* pin addr_2
* pin addr_3
* pin addr_4
* pin addr_5
* pin wl_7
* pin wl_8
* pin wl_9
* pin wl_10
* pin wl_11
* pin wl_12
* pin wl_13
* pin wl_14
* pin wl_15
* pin wl_16
* pin wl_17
* pin wl_18
* pin wl_19
* pin wl_20
* pin wl_21
* pin wl_22
* pin wl_23
* pin wl_24
* pin wl_25
* pin wl_26
* pin wl_27
* pin wl_28
* pin wl_29
* pin wl_30
* pin wl_31
* pin wl_32
* pin wl_33
* pin wl_34
* pin wl_35
* pin wl_36
* pin wl_37
* pin wl_38
* pin wl_39
* pin wl_40
* pin wl_41
* pin wl_42
* pin wl_43
* pin wl_44
* pin wl_45
* pin wl_46
* pin wl_47
* pin wl_48
* pin wl_49
* pin wl_50
* pin wl_51
* pin wl_52
* pin wl_53
* pin wl_54
* pin wl_55
* pin wl_56
* pin wl_57
* pin wl_58
* pin wl_59
* pin wl_60
* pin wl_61
* pin wl_62
* pin wl_63
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_port_address 1 2 5 7 9 10 13 14 17 18
+ 19 20 21 22 23 24 27 28 31 33 35 36 39 40 43 44 47 48 51 52 55 56 59 60 63 64
+ 67 68 71 72 75 76 79 80 83 84 87 88 91 92 95 96 99 100 103 104 107 108 111
+ 112 115 116 119 120 123 124 127 128 131 132 135 136 137 138
* net 1 wl_en
* net 2 rbl_wl
* net 5 wl_0
* net 7 wl_1
* net 9 wl_2
* net 10 wl_3
* net 13 wl_4
* net 14 wl_5
* net 17 wl_6
* net 18 addr_0
* net 19 addr_1
* net 20 addr_2
* net 21 addr_3
* net 22 addr_4
* net 23 addr_5
* net 24 wl_7
* net 27 wl_8
* net 28 wl_9
* net 31 wl_10
* net 33 wl_11
* net 35 wl_12
* net 36 wl_13
* net 39 wl_14
* net 40 wl_15
* net 43 wl_16
* net 44 wl_17
* net 47 wl_18
* net 48 wl_19
* net 51 wl_20
* net 52 wl_21
* net 55 wl_22
* net 56 wl_23
* net 59 wl_24
* net 60 wl_25
* net 63 wl_26
* net 64 wl_27
* net 67 wl_28
* net 68 wl_29
* net 71 wl_30
* net 72 wl_31
* net 75 wl_32
* net 76 wl_33
* net 79 wl_34
* net 80 wl_35
* net 83 wl_36
* net 84 wl_37
* net 87 wl_38
* net 88 wl_39
* net 91 wl_40
* net 92 wl_41
* net 95 wl_42
* net 96 wl_43
* net 99 wl_44
* net 100 wl_45
* net 103 wl_46
* net 104 wl_47
* net 107 wl_48
* net 108 wl_49
* net 111 wl_50
* net 112 wl_51
* net 115 wl_52
* net 116 wl_53
* net 119 wl_54
* net 120 wl_55
* net 123 wl_56
* net 124 wl_57
* net 127 wl_58
* net 128 wl_59
* net 131 wl_60
* net 132 wl_61
* net 135 wl_62
* net 136 wl_63
* net 137 vdd
* net 138 gnd
* cell instance $1 r0 *1 8.515,0
X$1 3 5 4 7 6 9 8 10 12 13 11 14 16 17 15 24 26 27 25 28 29 31 30 33 32 35 34
+ 36 37 39 38 40 42 43 41 44 46 47 45 48 50 51 49 52 54 55 53 56 58 59 57 60 62
+ 63 61 64 66 67 65 68 70 71 69 1 72 73 75 76 74 77 79 80 78 81 83 84 82 85 87
+ 88 86 89 91 92 90 93 95 96 94 97 99 100 98 101 103 104 102 105 107 108 106
+ 109 111 112 110 113 115 116 114 117 119 120 118 121 123 124 122 125 127 128
+ 126 129 131 132 130 133 135 136 134 137 138
+ custom_sram_1r1w_32_256_freepdk45_wordline_driver_array
* cell instance $2 m0 *1 9.075,0
X$2 1 2 137 138 custom_sram_1r1w_32_256_freepdk45_pinv_2
* cell instance $4 r0 *1 0,0
X$4 4 3 19 18 6 8 11 12 15 16 20 21 22 23 26 29 30 25 32 37 34 41 42 38 46 45
+ 50 49 54 53 58 57 62 61 66 65 70 69 73 74 77 78 81 82 85 86 89 90 93 94 97 98
+ 101 102 105 106 109 110 113 114 117 118 121 122 125 126 129 130 133 134 137
+ 138 custom_sram_1r1w_32_256_freepdk45_hierarchical_decoder
.ENDS custom_sram_1r1w_32_256_freepdk45_port_address

* cell custom_sram_1r1w_32_256_freepdk45_port_data_0
* pin bl_0
* pin br_0
* pin bl_1
* pin br_1
* pin bl_2
* pin bl_3
* pin bl_4
* pin br_4
* pin bl_5
* pin br_5
* pin bl_6
* pin br_6
* pin bl_7
* pin br_7
* pin bl_8
* pin br_8
* pin bl_9
* pin br_9
* pin bl_10
* pin br_10
* pin bl_11
* pin br_11
* pin bl_12
* pin br_12
* pin bl_13
* pin bl_14
* pin br_14
* pin bl_15
* pin br_15
* pin bl_16
* pin bl_17
* pin br_17
* pin bl_18
* pin br_18
* pin bl_19
* pin br_19
* pin bl_20
* pin br_20
* pin bl_21
* pin br_21
* pin bl_22
* pin br_22
* pin bl_23
* pin br_23
* pin bl_24
* pin br_24
* pin bl_25
* pin br_25
* pin bl_26
* pin br_26
* pin bl_27
* pin br_27
* pin bl_28
* pin br_28
* pin bl_29
* pin br_29
* pin bl_30
* pin br_30
* pin bl_31
* pin br_31
* pin bl_32
* pin br_32
* pin bl_33
* pin bl_34
* pin br_34
* pin bl_35
* pin bl_36
* pin br_36
* pin bl_37
* pin br_37
* pin bl_38
* pin br_38
* pin bl_39
* pin br_39
* pin bl_40
* pin br_40
* pin bl_41
* pin br_41
* pin bl_42
* pin br_42
* pin bl_43
* pin bl_44
* pin br_44
* pin bl_45
* pin bl_46
* pin br_46
* pin bl_47
* pin br_47
* pin bl_48
* pin br_48
* pin bl_49
* pin br_49
* pin bl_50
* pin br_50
* pin bl_51
* pin br_51
* pin bl_52
* pin bl_53
* pin br_53
* pin bl_54
* pin br_54
* pin bl_55
* pin br_55
* pin bl_56
* pin br_56
* pin bl_57
* pin br_57
* pin bl_58
* pin br_58
* pin bl_59
* pin br_59
* pin bl_60
* pin br_60
* pin bl_61
* pin br_61
* pin bl_62
* pin br_62
* pin bl_63
* pin br_63
* pin bl_64
* pin br_64
* pin bl_65
* pin br_65
* pin bl_66
* pin br_66
* pin bl_67
* pin br_67
* pin bl_68
* pin br_68
* pin bl_69
* pin br_69
* pin bl_70
* pin br_70
* pin bl_71
* pin bl_72
* pin br_72
* pin bl_73
* pin br_73
* pin bl_74
* pin br_74
* pin bl_75
* pin bl_76
* pin br_76
* pin bl_77
* pin br_77
* pin bl_78
* pin br_78
* pin bl_79
* pin br_79
* pin bl_80
* pin br_80
* pin bl_81
* pin bl_82
* pin bl_83
* pin br_83
* pin bl_84
* pin br_84
* pin bl_85
* pin br_85
* pin bl_86
* pin br_86
* pin bl_87
* pin br_87
* pin bl_88
* pin br_88
* pin bl_89
* pin br_89
* pin bl_90
* pin br_90
* pin bl_91
* pin br_91
* pin bl_92
* pin br_92
* pin bl_93
* pin br_93
* pin bl_94
* pin bl_95
* pin br_95
* pin bl_96
* pin br_96
* pin bl_97
* pin br_97
* pin bl_98
* pin br_98
* pin bl_99
* pin br_99
* pin bl_100
* pin br_100
* pin bl_101
* pin br_101
* pin bl_102
* pin br_102
* pin bl_103
* pin br_103
* pin bl_104
* pin br_104
* pin bl_105
* pin br_105
* pin bl_106
* pin br_106
* pin bl_107
* pin bl_108
* pin br_108
* pin bl_109
* pin bl_110
* pin br_110
* pin bl_111
* pin br_111
* pin bl_112
* pin br_112
* pin bl_113
* pin br_113
* pin bl_114
* pin br_114
* pin bl_115
* pin br_115
* pin bl_116
* pin br_116
* pin bl_117
* pin br_117
* pin bl_118
* pin br_118
* pin bl_119
* pin br_119
* pin bl_120
* pin br_120
* pin bl_121
* pin br_121
* pin bl_122
* pin br_122
* pin bl_123
* pin br_123
* pin bl_124
* pin br_124
* pin bl_125
* pin br_125
* pin bl_126
* pin br_126
* pin bl_127
* pin br_127
* pin rbl_bl
* pin rbl_br
* pin br_2
* pin br_3
* pin br_13
* pin br_16
* pin br_33
* pin br_35
* pin br_43
* pin br_45
* pin br_52
* pin p_en_bar
* pin br_71
* pin br_75
* pin br_81
* pin br_82
* pin br_94
* pin br_107
* pin br_109
* pin dout_0
* pin dout_1
* pin dout_2
* pin dout_3
* pin dout_4
* pin dout_5
* pin dout_6
* pin dout_7
* pin dout_8
* pin dout_9
* pin dout_10
* pin dout_11
* pin dout_12
* pin dout_13
* pin dout_14
* pin dout_15
* pin s_en
* pin sel_3
* pin sel_2
* pin sel_0
* pin sel_1
* pin dout_16
* pin dout_17
* pin dout_18
* pin dout_19
* pin dout_20
* pin dout_21
* pin dout_22
* pin dout_23
* pin dout_24
* pin dout_25
* pin dout_26
* pin dout_27
* pin dout_28
* pin dout_29
* pin dout_30
* pin dout_31
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_port_data_0 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37
+ 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89
+ 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111
+ 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130
+ 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149
+ 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168
+ 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187
+ 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206
+ 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225
+ 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244
+ 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 263 266 269
+ 272 275 278 281 284 287 290 293 296 299 302 305 308 309 310 311 312 313 316
+ 319 322 325 328 331 334 337 340 343 346 349 352 355 358 361 362
* net 1 bl_0
* net 2 br_0
* net 3 bl_1
* net 4 br_1
* net 5 bl_2
* net 6 bl_3
* net 7 bl_4
* net 8 br_4
* net 9 bl_5
* net 10 br_5
* net 11 bl_6
* net 12 br_6
* net 13 bl_7
* net 14 br_7
* net 15 bl_8
* net 16 br_8
* net 17 bl_9
* net 18 br_9
* net 19 bl_10
* net 20 br_10
* net 21 bl_11
* net 22 br_11
* net 23 bl_12
* net 24 br_12
* net 25 bl_13
* net 26 bl_14
* net 27 br_14
* net 28 bl_15
* net 29 br_15
* net 30 bl_16
* net 31 bl_17
* net 32 br_17
* net 33 bl_18
* net 34 br_18
* net 35 bl_19
* net 36 br_19
* net 37 bl_20
* net 38 br_20
* net 39 bl_21
* net 40 br_21
* net 41 bl_22
* net 42 br_22
* net 43 bl_23
* net 44 br_23
* net 45 bl_24
* net 46 br_24
* net 47 bl_25
* net 48 br_25
* net 49 bl_26
* net 50 br_26
* net 51 bl_27
* net 52 br_27
* net 53 bl_28
* net 54 br_28
* net 55 bl_29
* net 56 br_29
* net 57 bl_30
* net 58 br_30
* net 59 bl_31
* net 60 br_31
* net 61 bl_32
* net 62 br_32
* net 63 bl_33
* net 64 bl_34
* net 65 br_34
* net 66 bl_35
* net 67 bl_36
* net 68 br_36
* net 69 bl_37
* net 70 br_37
* net 71 bl_38
* net 72 br_38
* net 73 bl_39
* net 74 br_39
* net 75 bl_40
* net 76 br_40
* net 77 bl_41
* net 78 br_41
* net 79 bl_42
* net 80 br_42
* net 81 bl_43
* net 82 bl_44
* net 83 br_44
* net 84 bl_45
* net 85 bl_46
* net 86 br_46
* net 87 bl_47
* net 88 br_47
* net 89 bl_48
* net 90 br_48
* net 91 bl_49
* net 92 br_49
* net 93 bl_50
* net 94 br_50
* net 95 bl_51
* net 96 br_51
* net 97 bl_52
* net 98 bl_53
* net 99 br_53
* net 100 bl_54
* net 101 br_54
* net 102 bl_55
* net 103 br_55
* net 104 bl_56
* net 105 br_56
* net 106 bl_57
* net 107 br_57
* net 108 bl_58
* net 109 br_58
* net 110 bl_59
* net 111 br_59
* net 112 bl_60
* net 113 br_60
* net 114 bl_61
* net 115 br_61
* net 116 bl_62
* net 117 br_62
* net 118 bl_63
* net 119 br_63
* net 120 bl_64
* net 121 br_64
* net 122 bl_65
* net 123 br_65
* net 124 bl_66
* net 125 br_66
* net 126 bl_67
* net 127 br_67
* net 128 bl_68
* net 129 br_68
* net 130 bl_69
* net 131 br_69
* net 132 bl_70
* net 133 br_70
* net 134 bl_71
* net 135 bl_72
* net 136 br_72
* net 137 bl_73
* net 138 br_73
* net 139 bl_74
* net 140 br_74
* net 141 bl_75
* net 142 bl_76
* net 143 br_76
* net 144 bl_77
* net 145 br_77
* net 146 bl_78
* net 147 br_78
* net 148 bl_79
* net 149 br_79
* net 150 bl_80
* net 151 br_80
* net 152 bl_81
* net 153 bl_82
* net 154 bl_83
* net 155 br_83
* net 156 bl_84
* net 157 br_84
* net 158 bl_85
* net 159 br_85
* net 160 bl_86
* net 161 br_86
* net 162 bl_87
* net 163 br_87
* net 164 bl_88
* net 165 br_88
* net 166 bl_89
* net 167 br_89
* net 168 bl_90
* net 169 br_90
* net 170 bl_91
* net 171 br_91
* net 172 bl_92
* net 173 br_92
* net 174 bl_93
* net 175 br_93
* net 176 bl_94
* net 177 bl_95
* net 178 br_95
* net 179 bl_96
* net 180 br_96
* net 181 bl_97
* net 182 br_97
* net 183 bl_98
* net 184 br_98
* net 185 bl_99
* net 186 br_99
* net 187 bl_100
* net 188 br_100
* net 189 bl_101
* net 190 br_101
* net 191 bl_102
* net 192 br_102
* net 193 bl_103
* net 194 br_103
* net 195 bl_104
* net 196 br_104
* net 197 bl_105
* net 198 br_105
* net 199 bl_106
* net 200 br_106
* net 201 bl_107
* net 202 bl_108
* net 203 br_108
* net 204 bl_109
* net 205 bl_110
* net 206 br_110
* net 207 bl_111
* net 208 br_111
* net 209 bl_112
* net 210 br_112
* net 211 bl_113
* net 212 br_113
* net 213 bl_114
* net 214 br_114
* net 215 bl_115
* net 216 br_115
* net 217 bl_116
* net 218 br_116
* net 219 bl_117
* net 220 br_117
* net 221 bl_118
* net 222 br_118
* net 223 bl_119
* net 224 br_119
* net 225 bl_120
* net 226 br_120
* net 227 bl_121
* net 228 br_121
* net 229 bl_122
* net 230 br_122
* net 231 bl_123
* net 232 br_123
* net 233 bl_124
* net 234 br_124
* net 235 bl_125
* net 236 br_125
* net 237 bl_126
* net 238 br_126
* net 239 bl_127
* net 240 br_127
* net 241 rbl_bl
* net 242 rbl_br
* net 243 br_2
* net 244 br_3
* net 245 br_13
* net 246 br_16
* net 247 br_33
* net 248 br_35
* net 249 br_43
* net 250 br_45
* net 251 br_52
* net 252 p_en_bar
* net 253 br_71
* net 254 br_75
* net 255 br_81
* net 256 br_82
* net 257 br_94
* net 258 br_107
* net 259 br_109
* net 260 dout_0
* net 263 dout_1
* net 266 dout_2
* net 269 dout_3
* net 272 dout_4
* net 275 dout_5
* net 278 dout_6
* net 281 dout_7
* net 284 dout_8
* net 287 dout_9
* net 290 dout_10
* net 293 dout_11
* net 296 dout_12
* net 299 dout_13
* net 302 dout_14
* net 305 dout_15
* net 308 s_en
* net 309 sel_3
* net 310 sel_2
* net 311 sel_0
* net 312 sel_1
* net 313 dout_16
* net 316 dout_17
* net 319 dout_18
* net 322 dout_19
* net 325 dout_20
* net 328 dout_21
* net 331 dout_22
* net 334 dout_23
* net 337 dout_24
* net 340 dout_25
* net 343 dout_26
* net 346 dout_27
* net 349 dout_28
* net 352 dout_29
* net 355 dout_30
* net 358 dout_31
* net 361 vdd
* net 362 gnd
* cell instance $1 m0 *1 0,1.845
X$1 252 1 2 3 4 5 243 6 244 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 245 26 27 28 29 30 246 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47
+ 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 247 64 65 66 248 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80 81 249 82 83 84 250 85 86 87 88 89 90 91 92 93
+ 94 95 96 97 251 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113
+ 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132
+ 133 134 253 135 136 137 138 139 140 141 254 142 143 144 145 146 147 148 149
+ 150 151 152 255 153 256 154 155 156 157 158 159 160 161 162 163 164 165 166
+ 167 168 169 170 171 172 173 174 175 176 257 177 178 179 180 181 182 183 184
+ 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 258 202
+ 203 204 259 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239
+ 240 241 242 361 custom_sram_1r1w_32_256_freepdk45_precharge_array_0
* cell instance $2 m0 *1 0,5.06
X$2 360 357 354 351 348 345 342 339 262 336 333 330 327 324 321 318 315 307 265
+ 304 301 298 295 292 289 286 283 280 268 277 274 271 311 312 359 261 356 353
+ 350 347 264 344 341 338 267 335 332 329 326 270 323 320 317 273 314 306 303
+ 300 276 297 294 291 279 288 285 282 310 309 1 2 3 4 5 243 6 244 7 8 9 10 11
+ 12 13 14 15 16 17 18 19 20 21 22 23 24 25 245 26 27 28 29 30 246 31 32 33 34
+ 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 247 64 65 66 248 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 249 82
+ 83 84 250 85 86 87 88 89 90 91 92 93 94 95 96 97 251 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 253 135 136 137 138 139 140
+ 141 254 142 143 144 145 146 147 148 149 150 151 152 255 153 256 154 155 156
+ 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175
+ 176 257 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193
+ 194 195 196 197 198 199 200 201 258 202 203 204 259 205 206 207 208 209 210
+ 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229
+ 230 231 232 233 234 235 236 237 238 239 240 362
+ custom_sram_1r1w_32_256_freepdk45_column_mux_array_0
* cell instance $3 m0 *1 0,11.575
X$3 260 263 266 269 272 275 278 281 284 287 290 293 296 299 302 305 313 316 319
+ 322 325 328 331 334 337 340 343 346 349 352 355 358 261 308 262 264 265 267
+ 268 270 271 273 274 276 277 279 280 282 283 285 286 288 289 291 292 294 295
+ 297 298 300 301 303 304 306 307 314 315 317 318 320 321 323 324 326 327 329
+ 330 332 333 335 336 338 339 341 342 344 345 347 348 350 351 353 354 356 357
+ 359 360 361 362 custom_sram_1r1w_32_256_freepdk45_sense_amp_array
.ENDS custom_sram_1r1w_32_256_freepdk45_port_data_0

* cell custom_sram_1r1w_32_256_freepdk45_port_data
* pin rbl_bl
* pin rbl_br
* pin bl_0
* pin br_0
* pin bl_1
* pin br_1
* pin bl_2
* pin br_2
* pin bl_3
* pin bl_4
* pin br_4
* pin bl_5
* pin br_5
* pin bl_6
* pin br_6
* pin bl_7
* pin br_7
* pin bl_8
* pin bl_9
* pin br_9
* pin bl_10
* pin br_10
* pin bl_11
* pin br_11
* pin bl_12
* pin br_12
* pin bl_13
* pin br_13
* pin bl_14
* pin br_14
* pin bl_15
* pin br_15
* pin bl_16
* pin bl_17
* pin bl_18
* pin bl_19
* pin bl_20
* pin br_20
* pin bl_21
* pin br_21
* pin bl_22
* pin br_22
* pin bl_23
* pin br_23
* pin bl_24
* pin bl_25
* pin bl_26
* pin bl_27
* pin br_27
* pin bl_28
* pin br_28
* pin bl_29
* pin br_29
* pin bl_30
* pin br_30
* pin bl_31
* pin br_31
* pin bl_32
* pin br_32
* pin bl_33
* pin br_33
* pin bl_34
* pin br_34
* pin bl_35
* pin br_35
* pin bl_36
* pin br_36
* pin bl_37
* pin br_37
* pin bl_38
* pin br_38
* pin bl_39
* pin bl_40
* pin br_40
* pin bl_41
* pin br_41
* pin bl_42
* pin br_42
* pin bl_43
* pin br_43
* pin bl_44
* pin bl_45
* pin bl_46
* pin br_46
* pin bl_47
* pin br_47
* pin bl_48
* pin br_48
* pin bl_49
* pin br_49
* pin bl_50
* pin br_50
* pin bl_51
* pin br_51
* pin bl_52
* pin br_52
* pin bl_53
* pin br_53
* pin bl_54
* pin br_54
* pin bl_55
* pin br_55
* pin bl_56
* pin br_56
* pin bl_57
* pin br_57
* pin bl_58
* pin br_58
* pin bl_59
* pin br_59
* pin bl_60
* pin br_60
* pin bl_61
* pin br_61
* pin bl_62
* pin br_62
* pin bl_63
* pin bl_64
* pin br_64
* pin bl_65
* pin br_65
* pin bl_66
* pin br_66
* pin bl_67
* pin br_67
* pin bl_68
* pin bl_69
* pin br_69
* pin bl_70
* pin br_70
* pin bl_71
* pin br_71
* pin bl_72
* pin bl_73
* pin br_73
* pin bl_74
* pin bl_75
* pin br_75
* pin bl_76
* pin br_76
* pin bl_77
* pin br_77
* pin bl_78
* pin br_78
* pin bl_79
* pin br_79
* pin bl_80
* pin br_80
* pin bl_81
* pin br_81
* pin bl_82
* pin br_82
* pin bl_83
* pin bl_84
* pin br_84
* pin bl_85
* pin br_85
* pin bl_86
* pin br_86
* pin bl_87
* pin br_87
* pin bl_88
* pin br_88
* pin bl_89
* pin br_89
* pin bl_90
* pin br_90
* pin bl_91
* pin br_91
* pin bl_92
* pin br_92
* pin bl_93
* pin br_93
* pin bl_94
* pin br_94
* pin bl_95
* pin br_95
* pin bl_96
* pin br_96
* pin bl_97
* pin br_97
* pin bl_98
* pin br_98
* pin bl_99
* pin br_99
* pin bl_100
* pin br_100
* pin bl_101
* pin br_101
* pin bl_102
* pin br_102
* pin bl_103
* pin bl_104
* pin bl_105
* pin br_105
* pin bl_106
* pin br_106
* pin bl_107
* pin br_107
* pin bl_108
* pin br_108
* pin bl_109
* pin br_109
* pin bl_110
* pin br_110
* pin bl_111
* pin bl_112
* pin bl_113
* pin br_113
* pin bl_114
* pin br_114
* pin bl_115
* pin br_115
* pin bl_116
* pin bl_117
* pin bl_118
* pin br_118
* pin bl_119
* pin br_119
* pin bl_120
* pin br_120
* pin bl_121
* pin br_121
* pin bl_122
* pin br_122
* pin bl_123
* pin br_123
* pin bl_124
* pin br_124
* pin bl_125
* pin br_125
* pin bl_126
* pin br_126
* pin bl_127
* pin br_127
* pin br_3
* pin br_8
* pin br_16
* pin br_17
* pin br_18
* pin br_19
* pin br_24
* pin br_25
* pin br_26
* pin br_39
* pin br_44
* pin br_45
* pin br_63
* pin p_en_bar
* pin br_68
* pin br_72
* pin br_74
* pin br_83
* pin br_103
* pin br_104
* pin br_111
* pin br_112
* pin br_116
* pin br_117
* pin din_0
* pin din_1
* pin din_2
* pin din_3
* pin din_4
* pin din_5
* pin din_6
* pin din_7
* pin din_8
* pin din_9
* pin din_10
* pin din_11
* pin din_12
* pin din_13
* pin din_14
* pin din_15
* pin w_en
* pin sel_1
* pin sel_3
* pin sel_2
* pin sel_0
* pin din_16
* pin din_17
* pin din_18
* pin din_19
* pin din_20
* pin din_21
* pin din_22
* pin din_23
* pin din_24
* pin din_25
* pin din_26
* pin din_27
* pin din_28
* pin din_29
* pin din_30
* pin din_31
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_port_data 1 2 3 4 5 6 7 8 9 10 11 12
+ 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38
+ 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64
+ 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90
+ 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111
+ 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130
+ 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149
+ 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168
+ 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187
+ 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206
+ 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225
+ 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244
+ 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 261 264 267 270
+ 273 276 279 282 285 288 291 294 297 300 303 306 308 309 310 311 312 314 317
+ 320 323 326 329 332 335 338 341 344 347 350 353 356 359 361 362
* net 1 rbl_bl
* net 2 rbl_br
* net 3 bl_0
* net 4 br_0
* net 5 bl_1
* net 6 br_1
* net 7 bl_2
* net 8 br_2
* net 9 bl_3
* net 10 bl_4
* net 11 br_4
* net 12 bl_5
* net 13 br_5
* net 14 bl_6
* net 15 br_6
* net 16 bl_7
* net 17 br_7
* net 18 bl_8
* net 19 bl_9
* net 20 br_9
* net 21 bl_10
* net 22 br_10
* net 23 bl_11
* net 24 br_11
* net 25 bl_12
* net 26 br_12
* net 27 bl_13
* net 28 br_13
* net 29 bl_14
* net 30 br_14
* net 31 bl_15
* net 32 br_15
* net 33 bl_16
* net 34 bl_17
* net 35 bl_18
* net 36 bl_19
* net 37 bl_20
* net 38 br_20
* net 39 bl_21
* net 40 br_21
* net 41 bl_22
* net 42 br_22
* net 43 bl_23
* net 44 br_23
* net 45 bl_24
* net 46 bl_25
* net 47 bl_26
* net 48 bl_27
* net 49 br_27
* net 50 bl_28
* net 51 br_28
* net 52 bl_29
* net 53 br_29
* net 54 bl_30
* net 55 br_30
* net 56 bl_31
* net 57 br_31
* net 58 bl_32
* net 59 br_32
* net 60 bl_33
* net 61 br_33
* net 62 bl_34
* net 63 br_34
* net 64 bl_35
* net 65 br_35
* net 66 bl_36
* net 67 br_36
* net 68 bl_37
* net 69 br_37
* net 70 bl_38
* net 71 br_38
* net 72 bl_39
* net 73 bl_40
* net 74 br_40
* net 75 bl_41
* net 76 br_41
* net 77 bl_42
* net 78 br_42
* net 79 bl_43
* net 80 br_43
* net 81 bl_44
* net 82 bl_45
* net 83 bl_46
* net 84 br_46
* net 85 bl_47
* net 86 br_47
* net 87 bl_48
* net 88 br_48
* net 89 bl_49
* net 90 br_49
* net 91 bl_50
* net 92 br_50
* net 93 bl_51
* net 94 br_51
* net 95 bl_52
* net 96 br_52
* net 97 bl_53
* net 98 br_53
* net 99 bl_54
* net 100 br_54
* net 101 bl_55
* net 102 br_55
* net 103 bl_56
* net 104 br_56
* net 105 bl_57
* net 106 br_57
* net 107 bl_58
* net 108 br_58
* net 109 bl_59
* net 110 br_59
* net 111 bl_60
* net 112 br_60
* net 113 bl_61
* net 114 br_61
* net 115 bl_62
* net 116 br_62
* net 117 bl_63
* net 118 bl_64
* net 119 br_64
* net 120 bl_65
* net 121 br_65
* net 122 bl_66
* net 123 br_66
* net 124 bl_67
* net 125 br_67
* net 126 bl_68
* net 127 bl_69
* net 128 br_69
* net 129 bl_70
* net 130 br_70
* net 131 bl_71
* net 132 br_71
* net 133 bl_72
* net 134 bl_73
* net 135 br_73
* net 136 bl_74
* net 137 bl_75
* net 138 br_75
* net 139 bl_76
* net 140 br_76
* net 141 bl_77
* net 142 br_77
* net 143 bl_78
* net 144 br_78
* net 145 bl_79
* net 146 br_79
* net 147 bl_80
* net 148 br_80
* net 149 bl_81
* net 150 br_81
* net 151 bl_82
* net 152 br_82
* net 153 bl_83
* net 154 bl_84
* net 155 br_84
* net 156 bl_85
* net 157 br_85
* net 158 bl_86
* net 159 br_86
* net 160 bl_87
* net 161 br_87
* net 162 bl_88
* net 163 br_88
* net 164 bl_89
* net 165 br_89
* net 166 bl_90
* net 167 br_90
* net 168 bl_91
* net 169 br_91
* net 170 bl_92
* net 171 br_92
* net 172 bl_93
* net 173 br_93
* net 174 bl_94
* net 175 br_94
* net 176 bl_95
* net 177 br_95
* net 178 bl_96
* net 179 br_96
* net 180 bl_97
* net 181 br_97
* net 182 bl_98
* net 183 br_98
* net 184 bl_99
* net 185 br_99
* net 186 bl_100
* net 187 br_100
* net 188 bl_101
* net 189 br_101
* net 190 bl_102
* net 191 br_102
* net 192 bl_103
* net 193 bl_104
* net 194 bl_105
* net 195 br_105
* net 196 bl_106
* net 197 br_106
* net 198 bl_107
* net 199 br_107
* net 200 bl_108
* net 201 br_108
* net 202 bl_109
* net 203 br_109
* net 204 bl_110
* net 205 br_110
* net 206 bl_111
* net 207 bl_112
* net 208 bl_113
* net 209 br_113
* net 210 bl_114
* net 211 br_114
* net 212 bl_115
* net 213 br_115
* net 214 bl_116
* net 215 bl_117
* net 216 bl_118
* net 217 br_118
* net 218 bl_119
* net 219 br_119
* net 220 bl_120
* net 221 br_120
* net 222 bl_121
* net 223 br_121
* net 224 bl_122
* net 225 br_122
* net 226 bl_123
* net 227 br_123
* net 228 bl_124
* net 229 br_124
* net 230 bl_125
* net 231 br_125
* net 232 bl_126
* net 233 br_126
* net 234 bl_127
* net 235 br_127
* net 236 br_3
* net 237 br_8
* net 238 br_16
* net 239 br_17
* net 240 br_18
* net 241 br_19
* net 242 br_24
* net 243 br_25
* net 244 br_26
* net 245 br_39
* net 246 br_44
* net 247 br_45
* net 248 br_63
* net 249 p_en_bar
* net 250 br_68
* net 251 br_72
* net 252 br_74
* net 253 br_83
* net 254 br_103
* net 255 br_104
* net 256 br_111
* net 257 br_112
* net 258 br_116
* net 259 br_117
* net 261 din_0
* net 264 din_1
* net 267 din_2
* net 270 din_3
* net 273 din_4
* net 276 din_5
* net 279 din_6
* net 282 din_7
* net 285 din_8
* net 288 din_9
* net 291 din_10
* net 294 din_11
* net 297 din_12
* net 300 din_13
* net 303 din_14
* net 306 din_15
* net 308 w_en
* net 309 sel_1
* net 310 sel_3
* net 311 sel_2
* net 312 sel_0
* net 314 din_16
* net 317 din_17
* net 320 din_18
* net 323 din_19
* net 326 din_20
* net 329 din_21
* net 332 din_22
* net 335 din_23
* net 338 din_24
* net 341 din_25
* net 344 din_26
* net 347 din_27
* net 350 din_28
* net 353 din_29
* net 356 din_30
* net 359 din_31
* net 361 vdd
* net 362 gnd
* cell instance $1 m0 *1 0,1.845
X$1 249 1 2 3 4 5 6 7 8 9 236 10 11 12 13 14 15 16 17 18 237 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 238 34 239 35 240 36 241 37 38 39 40 41 42 43 44
+ 45 242 46 243 47 244 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66
+ 67 68 69 70 71 72 245 73 74 75 76 77 78 79 80 81 246 82 247 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 248 118 119 120 121 122 123 124 125 126 250 127
+ 128 129 130 131 132 133 251 134 135 136 252 137 138 139 140 141 142 143 144
+ 145 146 147 148 149 150 151 152 153 253 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 254 193 255 194 195 196 197 198
+ 199 200 201 202 203 204 205 206 256 207 257 208 209 210 211 212 213 214 258
+ 215 259 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232
+ 233 234 235 361 custom_sram_1r1w_32_256_freepdk45_precharge_array
* cell instance $2 m0 *1 0,5.06
X$2 360 357 354 351 348 345 342 339 262 336 333 330 327 324 321 318 315 307 265
+ 304 301 298 295 292 289 286 283 280 268 277 274 271 312 309 358 260 355 352
+ 349 346 263 343 340 337 266 334 331 328 325 269 322 319 316 272 313 305 302
+ 299 275 296 293 290 278 287 284 281 311 310 3 4 5 6 7 8 9 236 10 11 12 13 14
+ 15 16 17 18 237 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 238 34 239 35
+ 240 36 241 37 38 39 40 41 42 43 44 45 242 46 243 47 244 48 49 50 51 52 53 54
+ 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 245 73 74 75 76 77 78
+ 79 80 81 246 82 247 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 248 118
+ 119 120 121 122 123 124 125 126 250 127 128 129 130 131 132 133 251 134 135
+ 136 252 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153
+ 253 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171
+ 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190
+ 191 192 254 193 255 194 195 196 197 198 199 200 201 202 203 204 205 206 256
+ 207 257 208 209 210 211 212 213 214 258 215 259 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 362
+ custom_sram_1r1w_32_256_freepdk45_column_mux_array
* cell instance $3 m0 *1 0,9.74
X$3 261 264 267 270 273 276 279 282 285 288 291 294 297 300 303 306 314 317 320
+ 323 326 329 332 335 338 341 344 347 350 353 356 359 262 265 268 271 274 277
+ 280 283 286 289 292 295 298 301 304 307 308 315 318 321 324 327 330 333 336
+ 339 342 345 348 351 354 357 360 260 263 266 269 272 275 278 281 284 287 290
+ 293 296 299 302 305 313 316 319 322 325 328 331 334 337 340 343 346 349 352
+ 355 358 361 362 custom_sram_1r1w_32_256_freepdk45_write_driver_array
.ENDS custom_sram_1r1w_32_256_freepdk45_port_data

* cell custom_sram_1r1w_32_256_freepdk45_global_bitcell_array
* pin wl_0_10
* pin wl_0_11
* pin wl_0_12
* pin wl_0_13
* pin wl_0_14
* pin wl_0_15
* pin wl_0_16
* pin wl_0_2
* pin wl_0_1
* pin wl_0_3
* pin wl_0_4
* pin wl_0_9
* pin wl_0_5
* pin wl_0_6
* pin wl_0_7
* pin wl_0_8
* pin wl_0_0
* pin rbl_wl_0_0
* pin wl_0_31
* pin wl_0_30
* pin wl_0_29
* pin wl_0_28
* pin wl_0_27
* pin wl_0_26
* pin wl_0_17
* pin wl_0_18
* pin wl_0_19
* pin wl_0_20
* pin wl_0_21
* pin wl_0_22
* pin wl_0_23
* pin wl_0_24
* pin wl_0_25
* pin rbl_bl_0_0
* pin rbl_br_0_0
* pin bl_0_0
* pin bl_1_0
* pin br_1_0
* pin br_0_0
* pin bl_0_1
* pin bl_1_1
* pin br_1_1
* pin br_0_1
* pin bl_0_2
* pin bl_1_2
* pin br_1_2
* pin br_0_2
* pin bl_0_3
* pin bl_1_3
* pin br_1_3
* pin br_0_3
* pin bl_0_4
* pin bl_1_4
* pin br_1_4
* pin br_0_4
* pin bl_0_5
* pin bl_1_5
* pin br_1_5
* pin br_0_5
* pin bl_0_6
* pin bl_1_6
* pin br_1_6
* pin br_0_6
* pin bl_0_7
* pin bl_1_7
* pin br_1_7
* pin br_0_7
* pin bl_0_8
* pin bl_1_8
* pin br_1_8
* pin br_0_8
* pin bl_0_9
* pin bl_1_9
* pin br_1_9
* pin br_0_9
* pin bl_0_10
* pin bl_1_10
* pin br_1_10
* pin br_0_10
* pin bl_0_11
* pin bl_1_11
* pin br_1_11
* pin br_0_11
* pin bl_0_12
* pin bl_1_12
* pin br_1_12
* pin br_0_12
* pin bl_0_13
* pin bl_1_13
* pin br_1_13
* pin br_0_13
* pin bl_0_14
* pin bl_1_14
* pin br_1_14
* pin br_0_14
* pin bl_0_15
* pin bl_1_15
* pin br_1_15
* pin br_0_15
* pin bl_0_16
* pin bl_1_16
* pin br_1_16
* pin br_0_16
* pin bl_0_17
* pin bl_1_17
* pin br_1_17
* pin br_0_17
* pin bl_0_18
* pin bl_1_18
* pin br_1_18
* pin br_0_18
* pin bl_0_19
* pin bl_1_19
* pin br_1_19
* pin br_0_19
* pin bl_0_20
* pin bl_1_20
* pin br_1_20
* pin br_0_20
* pin bl_0_21
* pin bl_1_21
* pin br_1_21
* pin br_0_21
* pin bl_0_22
* pin bl_1_22
* pin br_1_22
* pin br_0_22
* pin bl_0_23
* pin bl_1_23
* pin br_1_23
* pin br_0_23
* pin bl_0_24
* pin bl_1_24
* pin br_1_24
* pin br_0_24
* pin bl_0_25
* pin bl_1_25
* pin br_1_25
* pin br_0_25
* pin bl_0_26
* pin bl_1_26
* pin br_1_26
* pin br_0_26
* pin bl_0_27
* pin bl_1_27
* pin br_1_27
* pin br_0_27
* pin bl_0_28
* pin bl_1_28
* pin br_1_28
* pin br_0_28
* pin bl_0_29
* pin bl_1_29
* pin br_1_29
* pin br_0_29
* pin bl_0_30
* pin bl_1_30
* pin br_1_30
* pin br_0_30
* pin bl_0_31
* pin bl_1_31
* pin br_1_31
* pin br_0_31
* pin wl_1_17
* pin wl_1_12
* pin wl_1_16
* pin wl_1_13
* pin wl_1_11
* pin wl_1_5
* pin wl_1_15
* pin wl_1_4
* pin wl_1_6
* pin wl_1_14
* pin wl_1_31
* pin wl_1_24
* pin wl_1_25
* pin wl_1_26
* pin wl_1_9
* pin wl_1_30
* pin wl_1_29
* pin wl_1_27
* pin wl_1_28
* pin wl_1_0
* pin wl_1_18
* pin wl_1_3
* pin wl_1_2
* pin wl_1_19
* pin wl_1_7
* pin wl_1_1
* pin wl_1_20
* pin wl_1_21
* pin wl_1_8
* pin wl_1_22
* pin wl_1_10
* pin wl_1_23
* pin bl_0_32
* pin bl_1_32
* pin br_1_32
* pin br_0_32
* pin bl_0_33
* pin bl_1_33
* pin br_1_33
* pin br_0_33
* pin bl_0_34
* pin bl_1_34
* pin br_1_34
* pin br_0_34
* pin bl_0_35
* pin bl_1_35
* pin br_1_35
* pin br_0_35
* pin bl_0_36
* pin bl_1_36
* pin br_1_36
* pin br_0_36
* pin bl_0_37
* pin bl_1_37
* pin br_1_37
* pin br_0_37
* pin bl_0_38
* pin bl_1_38
* pin br_1_38
* pin br_0_38
* pin bl_0_39
* pin bl_1_39
* pin br_1_39
* pin br_0_39
* pin bl_0_40
* pin bl_1_40
* pin br_1_40
* pin br_0_40
* pin bl_0_41
* pin bl_1_41
* pin br_1_41
* pin br_0_41
* pin bl_0_42
* pin bl_1_42
* pin br_1_42
* pin br_0_42
* pin bl_0_43
* pin bl_1_43
* pin br_1_43
* pin br_0_43
* pin bl_0_44
* pin bl_1_44
* pin br_1_44
* pin br_0_44
* pin bl_0_45
* pin bl_1_45
* pin br_1_45
* pin br_0_45
* pin bl_0_46
* pin bl_1_46
* pin br_1_46
* pin br_0_46
* pin bl_0_47
* pin bl_1_47
* pin br_1_47
* pin br_0_47
* pin bl_0_48
* pin bl_1_48
* pin br_1_48
* pin br_0_48
* pin bl_0_49
* pin bl_1_49
* pin br_1_49
* pin br_0_49
* pin bl_0_50
* pin bl_1_50
* pin br_1_50
* pin br_0_50
* pin bl_0_51
* pin bl_1_51
* pin br_1_51
* pin br_0_51
* pin bl_0_52
* pin bl_1_52
* pin br_1_52
* pin br_0_52
* pin bl_0_53
* pin bl_1_53
* pin br_1_53
* pin br_0_53
* pin bl_0_54
* pin bl_1_54
* pin br_1_54
* pin br_0_54
* pin bl_0_55
* pin bl_1_55
* pin br_1_55
* pin br_0_55
* pin bl_0_56
* pin bl_1_56
* pin br_1_56
* pin br_0_56
* pin bl_0_57
* pin bl_1_57
* pin br_1_57
* pin br_0_57
* pin bl_0_58
* pin bl_1_58
* pin br_1_58
* pin br_0_58
* pin bl_0_59
* pin bl_1_59
* pin br_1_59
* pin br_0_59
* pin bl_0_60
* pin bl_1_60
* pin br_1_60
* pin br_0_60
* pin bl_0_61
* pin bl_1_61
* pin br_1_61
* pin br_0_61
* pin bl_0_62
* pin bl_1_62
* pin br_1_62
* pin br_0_62
* pin bl_0_63
* pin bl_1_63
* pin br_1_63
* pin br_0_63
* pin bl_0_64
* pin bl_1_64
* pin br_1_64
* pin br_0_64
* pin bl_0_65
* pin bl_1_65
* pin br_1_65
* pin br_0_65
* pin bl_0_66
* pin bl_1_66
* pin br_1_66
* pin br_0_66
* pin bl_0_67
* pin bl_1_67
* pin br_1_67
* pin br_0_67
* pin bl_0_68
* pin bl_1_68
* pin br_1_68
* pin br_0_68
* pin bl_0_69
* pin bl_1_69
* pin br_1_69
* pin br_0_69
* pin bl_0_70
* pin bl_1_70
* pin br_1_70
* pin br_0_70
* pin bl_0_71
* pin bl_1_71
* pin br_1_71
* pin br_0_71
* pin bl_0_72
* pin bl_1_72
* pin br_1_72
* pin br_0_72
* pin bl_0_73
* pin bl_1_73
* pin br_1_73
* pin br_0_73
* pin bl_0_74
* pin bl_1_74
* pin br_1_74
* pin br_0_74
* pin bl_0_75
* pin bl_1_75
* pin br_1_75
* pin br_0_75
* pin bl_0_76
* pin bl_1_76
* pin br_1_76
* pin br_0_76
* pin bl_0_77
* pin bl_1_77
* pin br_1_77
* pin br_0_77
* pin bl_0_78
* pin bl_1_78
* pin br_1_78
* pin br_0_78
* pin bl_0_79
* pin bl_1_79
* pin br_1_79
* pin br_0_79
* pin bl_0_80
* pin bl_1_80
* pin br_1_80
* pin br_0_80
* pin bl_0_81
* pin bl_1_81
* pin br_1_81
* pin br_0_81
* pin bl_0_82
* pin bl_1_82
* pin br_1_82
* pin br_0_82
* pin bl_0_83
* pin bl_1_83
* pin br_1_83
* pin br_0_83
* pin bl_0_84
* pin bl_1_84
* pin br_1_84
* pin br_0_84
* pin bl_0_85
* pin bl_1_85
* pin br_1_85
* pin br_0_85
* pin bl_0_86
* pin bl_1_86
* pin br_1_86
* pin br_0_86
* pin bl_0_87
* pin bl_1_87
* pin br_1_87
* pin br_0_87
* pin bl_0_88
* pin bl_1_88
* pin br_1_88
* pin br_0_88
* pin bl_0_89
* pin bl_1_89
* pin br_1_89
* pin br_0_89
* pin bl_0_90
* pin bl_1_90
* pin br_1_90
* pin br_0_90
* pin bl_0_91
* pin bl_1_91
* pin br_1_91
* pin br_0_91
* pin bl_0_92
* pin bl_1_92
* pin br_1_92
* pin br_0_92
* pin bl_0_93
* pin bl_1_93
* pin br_1_93
* pin br_0_93
* pin bl_0_94
* pin bl_1_94
* pin br_1_94
* pin br_0_94
* pin bl_0_95
* pin bl_1_95
* pin br_1_95
* pin br_0_95
* pin bl_0_96
* pin bl_1_96
* pin br_1_96
* pin br_0_96
* pin bl_0_97
* pin bl_1_97
* pin br_1_97
* pin br_0_97
* pin bl_0_98
* pin bl_1_98
* pin br_1_98
* pin br_0_98
* pin bl_0_99
* pin bl_1_99
* pin br_1_99
* pin br_0_99
* pin bl_0_100
* pin bl_1_100
* pin br_1_100
* pin br_0_100
* pin bl_0_101
* pin bl_1_101
* pin br_1_101
* pin br_0_101
* pin bl_0_102
* pin bl_1_102
* pin br_1_102
* pin br_0_102
* pin bl_0_103
* pin bl_1_103
* pin br_1_103
* pin br_0_103
* pin bl_0_104
* pin bl_1_104
* pin br_1_104
* pin br_0_104
* pin bl_0_105
* pin bl_1_105
* pin br_1_105
* pin br_0_105
* pin bl_0_106
* pin bl_1_106
* pin br_1_106
* pin br_0_106
* pin bl_0_107
* pin bl_1_107
* pin br_1_107
* pin br_0_107
* pin bl_0_108
* pin bl_1_108
* pin br_1_108
* pin br_0_108
* pin bl_0_109
* pin bl_1_109
* pin br_1_109
* pin br_0_109
* pin bl_0_110
* pin bl_1_110
* pin br_1_110
* pin br_0_110
* pin bl_0_111
* pin bl_1_111
* pin br_1_111
* pin br_0_111
* pin bl_0_112
* pin bl_1_112
* pin br_1_112
* pin br_0_112
* pin bl_0_113
* pin bl_1_113
* pin br_1_113
* pin br_0_113
* pin bl_0_114
* pin bl_1_114
* pin br_1_114
* pin br_0_114
* pin bl_0_115
* pin bl_1_115
* pin br_1_115
* pin br_0_115
* pin bl_0_116
* pin bl_1_116
* pin br_1_116
* pin br_0_116
* pin bl_0_117
* pin bl_1_117
* pin br_1_117
* pin br_0_117
* pin bl_0_118
* pin bl_1_118
* pin br_1_118
* pin br_0_118
* pin bl_0_119
* pin bl_1_119
* pin br_1_119
* pin br_0_119
* pin bl_0_120
* pin bl_1_120
* pin br_1_120
* pin br_0_120
* pin bl_0_121
* pin bl_1_121
* pin br_1_121
* pin br_0_121
* pin bl_0_122
* pin bl_1_122
* pin br_1_122
* pin br_0_122
* pin bl_0_123
* pin bl_1_123
* pin br_1_123
* pin br_0_123
* pin bl_0_124
* pin bl_1_124
* pin br_1_124
* pin br_0_124
* pin bl_0_125
* pin bl_1_125
* pin br_1_125
* pin br_0_125
* pin bl_0_126
* pin bl_1_126
* pin br_1_126
* pin br_0_126
* pin bl_0_127
* pin bl_1_127
* pin br_1_127
* pin br_0_127
* pin rbl_bl_1_1
* pin rbl_br_1_1
* pin wl_0_51
* pin wl_0_35
* pin wl_0_52
* pin wl_0_36
* pin wl_0_53
* pin wl_0_42
* pin wl_0_41
* pin wl_0_37
* pin wl_0_54
* pin wl_0_40
* pin wl_0_55
* pin wl_0_46
* pin wl_0_47
* pin wl_0_45
* pin wl_0_32
* pin wl_0_48
* pin wl_0_44
* pin wl_0_38
* pin wl_0_49
* pin wl_0_33
* pin wl_0_43
* pin wl_0_50
* pin wl_0_34
* pin wl_0_39
* pin wl_0_63
* pin wl_0_62
* pin wl_0_61
* pin wl_0_60
* pin wl_0_59
* pin wl_0_58
* pin wl_0_56
* pin wl_0_57
* pin wl_1_63
* pin wl_1_62
* pin wl_1_60
* pin rbl_wl_1_1
* pin wl_1_61
* pin wl_1_44
* pin wl_1_43
* pin wl_1_42
* pin wl_1_41
* pin wl_1_40
* pin wl_1_39
* pin wl_1_38
* pin wl_1_37
* pin wl_1_36
* pin wl_1_35
* pin wl_1_34
* pin wl_1_33
* pin wl_1_32
* pin wl_1_59
* pin wl_1_58
* pin wl_1_57
* pin wl_1_56
* pin wl_1_55
* pin wl_1_54
* pin wl_1_53
* pin wl_1_52
* pin wl_1_51
* pin wl_1_50
* pin wl_1_49
* pin wl_1_48
* pin wl_1_47
* pin wl_1_46
* pin wl_1_45
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_global_bitcell_array 1 2 3 4 5 6 7 8
+ 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34
+ 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129
+ 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148
+ 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167
+ 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186
+ 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205
+ 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224
+ 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243
+ 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262
+ 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319
+ 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338
+ 339 340 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357
+ 358 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376
+ 377 378 379 380 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395
+ 396 397 398 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413 414
+ 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433
+ 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451 452
+ 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471
+ 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509
+ 510 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528
+ 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547
+ 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566
+ 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 583 584 586 587
+ 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606
+ 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625
+ 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643 644
+ 645 646 647 648 649 650 651 652
* net 1 wl_0_10
* net 2 wl_0_11
* net 3 wl_0_12
* net 4 wl_0_13
* net 5 wl_0_14
* net 6 wl_0_15
* net 7 wl_0_16
* net 8 wl_0_2
* net 9 wl_0_1
* net 10 wl_0_3
* net 11 wl_0_4
* net 12 wl_0_9
* net 13 wl_0_5
* net 14 wl_0_6
* net 15 wl_0_7
* net 16 wl_0_8
* net 17 wl_0_0
* net 18 rbl_wl_0_0
* net 19 wl_0_31
* net 20 wl_0_30
* net 21 wl_0_29
* net 22 wl_0_28
* net 23 wl_0_27
* net 24 wl_0_26
* net 25 wl_0_17
* net 26 wl_0_18
* net 27 wl_0_19
* net 28 wl_0_20
* net 29 wl_0_21
* net 30 wl_0_22
* net 31 wl_0_23
* net 32 wl_0_24
* net 33 wl_0_25
* net 34 rbl_bl_0_0
* net 35 rbl_bl_1_0
* net 36 rbl_br_1_0
* net 37 rbl_br_0_0
* net 38 bl_0_0
* net 39 bl_1_0
* net 40 br_1_0
* net 41 br_0_0
* net 42 bl_0_1
* net 43 bl_1_1
* net 44 br_1_1
* net 45 br_0_1
* net 46 bl_0_2
* net 47 bl_1_2
* net 48 br_1_2
* net 49 br_0_2
* net 50 bl_0_3
* net 51 bl_1_3
* net 52 br_1_3
* net 53 br_0_3
* net 54 bl_0_4
* net 55 bl_1_4
* net 56 br_1_4
* net 57 br_0_4
* net 58 bl_0_5
* net 59 bl_1_5
* net 60 br_1_5
* net 61 br_0_5
* net 62 bl_0_6
* net 63 bl_1_6
* net 64 br_1_6
* net 65 br_0_6
* net 66 bl_0_7
* net 67 bl_1_7
* net 68 br_1_7
* net 69 br_0_7
* net 70 bl_0_8
* net 71 bl_1_8
* net 72 br_1_8
* net 73 br_0_8
* net 74 bl_0_9
* net 75 bl_1_9
* net 76 br_1_9
* net 77 br_0_9
* net 78 bl_0_10
* net 79 bl_1_10
* net 80 br_1_10
* net 81 br_0_10
* net 82 bl_0_11
* net 83 bl_1_11
* net 84 br_1_11
* net 85 br_0_11
* net 86 bl_0_12
* net 87 bl_1_12
* net 88 br_1_12
* net 89 br_0_12
* net 90 bl_0_13
* net 91 bl_1_13
* net 92 br_1_13
* net 93 br_0_13
* net 94 bl_0_14
* net 95 bl_1_14
* net 96 br_1_14
* net 97 br_0_14
* net 98 bl_0_15
* net 99 bl_1_15
* net 100 br_1_15
* net 101 br_0_15
* net 102 bl_0_16
* net 103 bl_1_16
* net 104 br_1_16
* net 105 br_0_16
* net 106 bl_0_17
* net 107 bl_1_17
* net 108 br_1_17
* net 109 br_0_17
* net 110 bl_0_18
* net 111 bl_1_18
* net 112 br_1_18
* net 113 br_0_18
* net 114 bl_0_19
* net 115 bl_1_19
* net 116 br_1_19
* net 117 br_0_19
* net 118 bl_0_20
* net 119 bl_1_20
* net 120 br_1_20
* net 121 br_0_20
* net 122 bl_0_21
* net 123 bl_1_21
* net 124 br_1_21
* net 125 br_0_21
* net 126 bl_0_22
* net 127 bl_1_22
* net 128 br_1_22
* net 129 br_0_22
* net 130 bl_0_23
* net 131 bl_1_23
* net 132 br_1_23
* net 133 br_0_23
* net 134 bl_0_24
* net 135 bl_1_24
* net 136 br_1_24
* net 137 br_0_24
* net 138 bl_0_25
* net 139 bl_1_25
* net 140 br_1_25
* net 141 br_0_25
* net 142 bl_0_26
* net 143 bl_1_26
* net 144 br_1_26
* net 145 br_0_26
* net 146 bl_0_27
* net 147 bl_1_27
* net 148 br_1_27
* net 149 br_0_27
* net 150 bl_0_28
* net 151 bl_1_28
* net 152 br_1_28
* net 153 br_0_28
* net 154 bl_0_29
* net 155 bl_1_29
* net 156 br_1_29
* net 157 br_0_29
* net 158 bl_0_30
* net 159 bl_1_30
* net 160 br_1_30
* net 161 br_0_30
* net 162 bl_0_31
* net 163 bl_1_31
* net 164 br_1_31
* net 165 br_0_31
* net 166 wl_1_17
* net 167 wl_1_12
* net 168 wl_1_16
* net 169 wl_1_13
* net 170 wl_1_11
* net 171 wl_1_5
* net 172 wl_1_15
* net 173 wl_1_4
* net 174 wl_1_6
* net 175 wl_1_14
* net 176 wl_1_31
* net 177 wl_1_24
* net 178 wl_1_25
* net 179 wl_1_26
* net 180 wl_1_9
* net 181 wl_1_30
* net 182 wl_1_29
* net 183 wl_1_27
* net 184 wl_1_28
* net 185 wl_1_0
* net 186 wl_1_18
* net 187 wl_1_3
* net 188 wl_1_2
* net 189 wl_1_19
* net 190 wl_1_7
* net 191 wl_1_1
* net 192 wl_1_20
* net 193 wl_1_21
* net 194 wl_1_8
* net 195 wl_1_22
* net 196 wl_1_10
* net 197 wl_1_23
* net 198 bl_0_32
* net 199 bl_1_32
* net 200 br_1_32
* net 201 br_0_32
* net 202 bl_0_33
* net 203 bl_1_33
* net 204 br_1_33
* net 205 br_0_33
* net 206 bl_0_34
* net 207 bl_1_34
* net 208 br_1_34
* net 209 br_0_34
* net 210 bl_0_35
* net 211 bl_1_35
* net 212 br_1_35
* net 213 br_0_35
* net 214 bl_0_36
* net 215 bl_1_36
* net 216 br_1_36
* net 217 br_0_36
* net 218 bl_0_37
* net 219 bl_1_37
* net 220 br_1_37
* net 221 br_0_37
* net 222 bl_0_38
* net 223 bl_1_38
* net 224 br_1_38
* net 225 br_0_38
* net 226 bl_0_39
* net 227 bl_1_39
* net 228 br_1_39
* net 229 br_0_39
* net 230 bl_0_40
* net 231 bl_1_40
* net 232 br_1_40
* net 233 br_0_40
* net 234 bl_0_41
* net 235 bl_1_41
* net 236 br_1_41
* net 237 br_0_41
* net 238 bl_0_42
* net 239 bl_1_42
* net 240 br_1_42
* net 241 br_0_42
* net 242 bl_0_43
* net 243 bl_1_43
* net 244 br_1_43
* net 245 br_0_43
* net 246 bl_0_44
* net 247 bl_1_44
* net 248 br_1_44
* net 249 br_0_44
* net 250 bl_0_45
* net 251 bl_1_45
* net 252 br_1_45
* net 253 br_0_45
* net 254 bl_0_46
* net 255 bl_1_46
* net 256 br_1_46
* net 257 br_0_46
* net 258 bl_0_47
* net 259 bl_1_47
* net 260 br_1_47
* net 261 br_0_47
* net 262 bl_0_48
* net 263 bl_1_48
* net 264 br_1_48
* net 265 br_0_48
* net 266 bl_0_49
* net 267 bl_1_49
* net 268 br_1_49
* net 269 br_0_49
* net 270 bl_0_50
* net 271 bl_1_50
* net 272 br_1_50
* net 273 br_0_50
* net 274 bl_0_51
* net 275 bl_1_51
* net 276 br_1_51
* net 277 br_0_51
* net 278 bl_0_52
* net 279 bl_1_52
* net 280 br_1_52
* net 281 br_0_52
* net 282 bl_0_53
* net 283 bl_1_53
* net 284 br_1_53
* net 285 br_0_53
* net 286 bl_0_54
* net 287 bl_1_54
* net 288 br_1_54
* net 289 br_0_54
* net 290 bl_0_55
* net 291 bl_1_55
* net 292 br_1_55
* net 293 br_0_55
* net 294 bl_0_56
* net 295 bl_1_56
* net 296 br_1_56
* net 297 br_0_56
* net 298 bl_0_57
* net 299 bl_1_57
* net 300 br_1_57
* net 301 br_0_57
* net 302 bl_0_58
* net 303 bl_1_58
* net 304 br_1_58
* net 305 br_0_58
* net 306 bl_0_59
* net 307 bl_1_59
* net 308 br_1_59
* net 309 br_0_59
* net 310 bl_0_60
* net 311 bl_1_60
* net 312 br_1_60
* net 313 br_0_60
* net 314 bl_0_61
* net 315 bl_1_61
* net 316 br_1_61
* net 317 br_0_61
* net 318 bl_0_62
* net 319 bl_1_62
* net 320 br_1_62
* net 321 br_0_62
* net 322 bl_0_63
* net 323 bl_1_63
* net 324 br_1_63
* net 325 br_0_63
* net 326 bl_0_64
* net 327 bl_1_64
* net 328 br_1_64
* net 329 br_0_64
* net 330 bl_0_65
* net 331 bl_1_65
* net 332 br_1_65
* net 333 br_0_65
* net 334 bl_0_66
* net 335 bl_1_66
* net 336 br_1_66
* net 337 br_0_66
* net 338 bl_0_67
* net 339 bl_1_67
* net 340 br_1_67
* net 341 br_0_67
* net 342 bl_0_68
* net 343 bl_1_68
* net 344 br_1_68
* net 345 br_0_68
* net 346 bl_0_69
* net 347 bl_1_69
* net 348 br_1_69
* net 349 br_0_69
* net 350 bl_0_70
* net 351 bl_1_70
* net 352 br_1_70
* net 353 br_0_70
* net 354 bl_0_71
* net 355 bl_1_71
* net 356 br_1_71
* net 357 br_0_71
* net 358 bl_0_72
* net 359 bl_1_72
* net 360 br_1_72
* net 361 br_0_72
* net 362 bl_0_73
* net 363 bl_1_73
* net 364 br_1_73
* net 365 br_0_73
* net 366 bl_0_74
* net 367 bl_1_74
* net 368 br_1_74
* net 369 br_0_74
* net 370 bl_0_75
* net 371 bl_1_75
* net 372 br_1_75
* net 373 br_0_75
* net 374 bl_0_76
* net 375 bl_1_76
* net 376 br_1_76
* net 377 br_0_76
* net 378 bl_0_77
* net 379 bl_1_77
* net 380 br_1_77
* net 381 br_0_77
* net 382 bl_0_78
* net 383 bl_1_78
* net 384 br_1_78
* net 385 br_0_78
* net 386 bl_0_79
* net 387 bl_1_79
* net 388 br_1_79
* net 389 br_0_79
* net 390 bl_0_80
* net 391 bl_1_80
* net 392 br_1_80
* net 393 br_0_80
* net 394 bl_0_81
* net 395 bl_1_81
* net 396 br_1_81
* net 397 br_0_81
* net 398 bl_0_82
* net 399 bl_1_82
* net 400 br_1_82
* net 401 br_0_82
* net 402 bl_0_83
* net 403 bl_1_83
* net 404 br_1_83
* net 405 br_0_83
* net 406 bl_0_84
* net 407 bl_1_84
* net 408 br_1_84
* net 409 br_0_84
* net 410 bl_0_85
* net 411 bl_1_85
* net 412 br_1_85
* net 413 br_0_85
* net 414 bl_0_86
* net 415 bl_1_86
* net 416 br_1_86
* net 417 br_0_86
* net 418 bl_0_87
* net 419 bl_1_87
* net 420 br_1_87
* net 421 br_0_87
* net 422 bl_0_88
* net 423 bl_1_88
* net 424 br_1_88
* net 425 br_0_88
* net 426 bl_0_89
* net 427 bl_1_89
* net 428 br_1_89
* net 429 br_0_89
* net 430 bl_0_90
* net 431 bl_1_90
* net 432 br_1_90
* net 433 br_0_90
* net 434 bl_0_91
* net 435 bl_1_91
* net 436 br_1_91
* net 437 br_0_91
* net 438 bl_0_92
* net 439 bl_1_92
* net 440 br_1_92
* net 441 br_0_92
* net 442 bl_0_93
* net 443 bl_1_93
* net 444 br_1_93
* net 445 br_0_93
* net 446 bl_0_94
* net 447 bl_1_94
* net 448 br_1_94
* net 449 br_0_94
* net 450 bl_0_95
* net 451 bl_1_95
* net 452 br_1_95
* net 453 br_0_95
* net 454 bl_0_96
* net 455 bl_1_96
* net 456 br_1_96
* net 457 br_0_96
* net 458 bl_0_97
* net 459 bl_1_97
* net 460 br_1_97
* net 461 br_0_97
* net 462 bl_0_98
* net 463 bl_1_98
* net 464 br_1_98
* net 465 br_0_98
* net 466 bl_0_99
* net 467 bl_1_99
* net 468 br_1_99
* net 469 br_0_99
* net 470 bl_0_100
* net 471 bl_1_100
* net 472 br_1_100
* net 473 br_0_100
* net 474 bl_0_101
* net 475 bl_1_101
* net 476 br_1_101
* net 477 br_0_101
* net 478 bl_0_102
* net 479 bl_1_102
* net 480 br_1_102
* net 481 br_0_102
* net 482 bl_0_103
* net 483 bl_1_103
* net 484 br_1_103
* net 485 br_0_103
* net 486 bl_0_104
* net 487 bl_1_104
* net 488 br_1_104
* net 489 br_0_104
* net 490 bl_0_105
* net 491 bl_1_105
* net 492 br_1_105
* net 493 br_0_105
* net 494 bl_0_106
* net 495 bl_1_106
* net 496 br_1_106
* net 497 br_0_106
* net 498 bl_0_107
* net 499 bl_1_107
* net 500 br_1_107
* net 501 br_0_107
* net 502 bl_0_108
* net 503 bl_1_108
* net 504 br_1_108
* net 505 br_0_108
* net 506 bl_0_109
* net 507 bl_1_109
* net 508 br_1_109
* net 509 br_0_109
* net 510 bl_0_110
* net 511 bl_1_110
* net 512 br_1_110
* net 513 br_0_110
* net 514 bl_0_111
* net 515 bl_1_111
* net 516 br_1_111
* net 517 br_0_111
* net 518 bl_0_112
* net 519 bl_1_112
* net 520 br_1_112
* net 521 br_0_112
* net 522 bl_0_113
* net 523 bl_1_113
* net 524 br_1_113
* net 525 br_0_113
* net 526 bl_0_114
* net 527 bl_1_114
* net 528 br_1_114
* net 529 br_0_114
* net 530 bl_0_115
* net 531 bl_1_115
* net 532 br_1_115
* net 533 br_0_115
* net 534 bl_0_116
* net 535 bl_1_116
* net 536 br_1_116
* net 537 br_0_116
* net 538 bl_0_117
* net 539 bl_1_117
* net 540 br_1_117
* net 541 br_0_117
* net 542 bl_0_118
* net 543 bl_1_118
* net 544 br_1_118
* net 545 br_0_118
* net 546 bl_0_119
* net 547 bl_1_119
* net 548 br_1_119
* net 549 br_0_119
* net 550 bl_0_120
* net 551 bl_1_120
* net 552 br_1_120
* net 553 br_0_120
* net 554 bl_0_121
* net 555 bl_1_121
* net 556 br_1_121
* net 557 br_0_121
* net 558 bl_0_122
* net 559 bl_1_122
* net 560 br_1_122
* net 561 br_0_122
* net 562 bl_0_123
* net 563 bl_1_123
* net 564 br_1_123
* net 565 br_0_123
* net 566 bl_0_124
* net 567 bl_1_124
* net 568 br_1_124
* net 569 br_0_124
* net 570 bl_0_125
* net 571 bl_1_125
* net 572 br_1_125
* net 573 br_0_125
* net 574 bl_0_126
* net 575 bl_1_126
* net 576 br_1_126
* net 577 br_0_126
* net 578 bl_0_127
* net 579 bl_1_127
* net 580 br_1_127
* net 581 br_0_127
* net 582 rbl_bl_0_1
* net 583 rbl_bl_1_1
* net 584 rbl_br_1_1
* net 585 rbl_br_0_1
* net 586 wl_0_51
* net 587 wl_0_35
* net 588 wl_0_52
* net 589 wl_0_36
* net 590 wl_0_53
* net 591 wl_0_42
* net 592 wl_0_41
* net 593 wl_0_37
* net 594 wl_0_54
* net 595 wl_0_40
* net 596 wl_0_55
* net 597 wl_0_46
* net 598 wl_0_47
* net 599 wl_0_45
* net 600 wl_0_32
* net 601 wl_0_48
* net 602 wl_0_44
* net 603 wl_0_38
* net 604 wl_0_49
* net 605 wl_0_33
* net 606 wl_0_43
* net 607 wl_0_50
* net 608 wl_0_34
* net 609 wl_0_39
* net 610 wl_0_63
* net 611 wl_0_62
* net 612 wl_0_61
* net 613 wl_0_60
* net 614 wl_0_59
* net 615 wl_0_58
* net 616 wl_0_56
* net 617 wl_0_57
* net 618 wl_1_63
* net 619 wl_1_62
* net 620 wl_1_60
* net 621 rbl_wl_1_1
* net 622 wl_1_61
* net 623 wl_1_44
* net 624 wl_1_43
* net 625 wl_1_42
* net 626 wl_1_41
* net 627 wl_1_40
* net 628 wl_1_39
* net 629 wl_1_38
* net 630 wl_1_37
* net 631 wl_1_36
* net 632 wl_1_35
* net 633 wl_1_34
* net 634 wl_1_33
* net 635 wl_1_32
* net 636 wl_1_59
* net 637 wl_1_58
* net 638 wl_1_57
* net 639 wl_1_56
* net 640 wl_1_55
* net 641 wl_1_54
* net 642 wl_1_53
* net 643 wl_1_52
* net 644 wl_1_51
* net 645 wl_1_50
* net 646 wl_1_49
* net 647 wl_1_48
* net 648 wl_1_47
* net 649 wl_1_46
* net 650 wl_1_45
* net 651 vdd
* net 652 gnd
* cell instance $1 r0 *1 0,0
X$1 10 11 18 9 17 14 8 13 191 185 174 188 173 187 171 12 1 16 2 3 15 4 5 190
+ 169 194 180 196 170 167 28 25 7 26 27 6 29 172 175 193 186 189 166 168 192 23
+ 32 22 31 21 30 24 33 177 195 183 184 178 179 197 20 19 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66
+ 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92
+ 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113
+ 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132
+ 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151
+ 152 153 154 155 156 157 158 159 160 161 162 163 164 165 182 181 176 602 606
+ 593 603 591 609 592 595 600 605 597 599 589 587 608 623 649 633 634 632 650
+ 625 629 628 635 626 627 631 630 624 594 604 588 598 601 590 586 607 642 648
+ 645 644 646 643 647 614 613 596 615 612 617 611 616 641 639 636 622 620 637
+ 638 640 610 621 618 619 651 652
+ custom_sram_1r1w_32_256_freepdk45_local_bitcell_array
* cell instance $2 r0 *1 56.08,0
X$2 9 8 10 11 17 18 14 13 171 191 187 185 188 173 4 12 3 1 16 15 2 174 190 169
+ 196 170 180 194 167 25 26 7 6 27 29 5 28 172 192 175 189 168 166 186 32 31 33
+ 24 30 23 22 184 183 193 177 178 197 179 195 20 21 19 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279
+ 280 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298
+ 299 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317
+ 318 319 320 321 322 323 324 325 176 182 181 593 608 603 609 587 595 591 592
+ 600 605 589 597 599 606 602 633 627 650 628 629 632 635 634 624 625 630 623
+ 631 626 590 598 588 601 586 607 604 647 642 644 649 645 643 648 646 617 615
+ 596 616 614 613 612 594 640 620 641 636 639 638 637 611 610 621 622 618 619
+ 651 652 custom_sram_1r1w_32_256_freepdk45_local_bitcell_array_0
* cell instance $3 r0 *1 165.89,0
X$3 10 11 18 9 17 14 8 13 191 185 174 188 173 187 171 12 1 16 2 3 15 4 5 190
+ 169 194 180 196 170 167 28 25 7 26 27 6 29 172 175 193 186 189 166 168 192 23
+ 32 22 31 21 30 24 33 177 195 183 184 178 179 197 20 19 454 455 456 457 458
+ 459 460 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477
+ 478 479 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496
+ 497 498 499 500 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515
+ 516 517 518 519 520 521 522 523 524 525 526 527 528 529 530 531 532 533 534
+ 535 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550 551 552 553
+ 554 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570 571 572
+ 573 574 575 576 577 578 579 580 581 582 583 584 585 182 181 176 602 606 593
+ 603 591 609 592 595 600 605 597 599 589 587 608 623 649 633 634 632 650 625
+ 629 628 635 626 627 631 630 624 594 604 588 598 601 590 586 607 642 648 645
+ 644 646 643 647 614 613 596 615 612 617 611 616 641 639 636 622 620 637 638
+ 640 610 621 618 619 651 652
+ custom_sram_1r1w_32_256_freepdk45_local_bitcell_array_1
* cell instance $4 r0 *1 110.985,0
X$4 9 8 10 11 17 18 14 13 171 191 187 185 188 173 4 12 3 1 16 15 2 174 190 169
+ 196 170 180 194 167 25 26 7 6 27 29 5 28 172 192 175 189 168 166 186 32 31 33
+ 24 30 23 22 184 183 193 177 178 197 179 195 20 21 19 326 327 328 329 330 331
+ 332 333 334 335 336 337 338 339 340 341 342 343 344 345 346 347 348 349 350
+ 351 352 353 354 355 356 357 358 359 360 361 362 363 364 365 366 367 368 369
+ 370 371 372 373 374 375 376 377 378 379 380 381 382 383 384 385 386 387 388
+ 389 390 391 392 393 394 395 396 397 398 399 400 401 402 403 404 405 406 407
+ 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426
+ 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445
+ 446 447 448 449 450 451 452 453 176 182 181 593 608 603 609 587 595 591 592
+ 600 605 589 597 599 606 602 633 627 650 628 629 632 635 634 624 625 630 623
+ 631 626 590 598 588 601 586 607 604 647 642 644 649 645 643 648 646 617 615
+ 596 616 614 613 612 594 640 620 641 636 639 638 637 611 610 621 622 618 619
+ 651 652 custom_sram_1r1w_32_256_freepdk45_local_bitcell_array_0
.ENDS custom_sram_1r1w_32_256_freepdk45_global_bitcell_array

* cell custom_sram_1r1w_32_256_freepdk45_pdriver_3
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pdriver_3 1 2 3 4
* net 1 Z
* net 2 A
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 custom_sram_1r1w_32_256_freepdk45_pinv_16
.ENDS custom_sram_1r1w_32_256_freepdk45_pdriver_3

* cell custom_sram_1r1w_32_256_freepdk45_pinv_21
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_21 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.2735 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=3.8675U AS=0.43955625P AD=0.43955625P PS=7.12U
+ PD=7.12U
* device instance $14 r0 *1 0.2325,1.8985 PMOS_VTG
M$14 3 1 2 3 PMOS_VTG L=0.05U W=11.6025U AS=1.31866875P AD=1.31866875P
+ PS=15.45U PD=15.45U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_21

* cell custom_sram_1r1w_32_256_freepdk45_pinv_20
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_20 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.251 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=1.2625U AS=0.14581875P AD=0.14581875P PS=2.67U
+ PD=2.67U
* device instance $6 r0 *1 0.2325,1.9675 PMOS_VTG
M$6 3 1 2 3 PMOS_VTG L=0.05U W=3.775U AS=0.4360125P AD=0.4360125P PS=5.685U
+ PD=5.685U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_20

* cell custom_sram_1r1w_32_256_freepdk45_pinv_19
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_19 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.2375 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.45U AS=0.054P AD=0.054P PS=1.155U PD=1.155U
* device instance $3 r0 *1 0.2325,2.0075 PMOS_VTG
M$3 3 1 2 3 PMOS_VTG L=0.05U W=1.35U AS=0.162P AD=0.162P PS=2.505U PD=2.505U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_19

* cell custom_sram_1r1w_32_256_freepdk45_pinv_18
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_18 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.215 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.02295P PS=0.615U PD=0.615U
* device instance $2 r0 *1 0.2325,2.075 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.54U AS=0.06885P AD=0.06885P PS=1.335U PD=1.335U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_18

* cell custom_sram_1r1w_32_256_freepdk45_pinv_22
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_22 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.17 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.09U AS=0.011475P AD=0.011475P PS=0.435U
+ PD=0.435U
* device instance $2 r0 *1 0.2325,2.21 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_22

* cell custom_sram_1r1w_32_256_freepdk45_pdriver_4
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pdriver_4 1 2 3 4
* net 1 Z
* net 2 A
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 custom_sram_1r1w_32_256_freepdk45_pinv_17
.ENDS custom_sram_1r1w_32_256_freepdk45_pdriver_4

* cell custom_sram_1r1w_32_256_freepdk45_pnand3_0
* pin A
* pin B
* pin C
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pnand3_0 1 2 3 4 5 6
* net 1 A
* net 2 B
* net 3 C
* net 4 Z
* net 5 vdd
* net 6 gnd
* device instance $1 r0 *1 0.2325,2.21 PMOS_VTG
M$1 5 1 4 5 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,2.21 PMOS_VTG
M$2 4 2 5 5 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.022275P PS=0.435U
+ PD=0.435U
* device instance $3 r0 *1 0.6625,2.21 PMOS_VTG
M$3 5 3 4 5 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $4 r0 *1 0.2325,0.215 NMOS_VTG
M$4 6 1 8 6 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $5 r0 *1 0.4475,0.215 NMOS_VTG
M$5 8 2 7 6 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.01485P PS=0.345U PD=0.345U
* device instance $6 r0 *1 0.6625,0.215 NMOS_VTG
M$6 7 3 4 6 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS custom_sram_1r1w_32_256_freepdk45_pnand3_0

* cell custom_sram_1r1w_32_256_freepdk45_pinv_15
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_15 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.26 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=1.89U AS=0.216675P AD=0.216675P PS=3.765U
+ PD=3.765U
* device instance $8 r0 *1 0.2325,1.94 PMOS_VTG
M$8 3 1 2 3 PMOS_VTG L=0.05U W=5.67U AS=0.650025P AD=0.650025P PS=8.085U
+ PD=8.085U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_15

* cell custom_sram_1r1w_32_256_freepdk45_pinv_14
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_14 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.23 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.63U AS=0.074025P AD=0.074025P PS=1.545U
+ PD=1.545U
* device instance $4 r0 *1 0.2325,2.03 PMOS_VTG
M$4 3 1 2 3 PMOS_VTG L=0.05U W=1.89U AS=0.222075P AD=0.222075P PS=3.225U
+ PD=3.225U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_14

* cell custom_sram_1r1w_32_256_freepdk45_pdriver_0
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pdriver_0 1 2 3 4
* net 1 Z
* net 2 A
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 custom_sram_1r1w_32_256_freepdk45_pinv_7
.ENDS custom_sram_1r1w_32_256_freepdk45_pdriver_0

* cell custom_sram_1r1w_32_256_freepdk45_pinv_13
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_13 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.2735 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=6.545U AS=0.740775P AD=0.740775P PS=11.8225U
+ PD=11.8225U
* device instance $23 r0 *1 0.2325,1.8975 PMOS_VTG
M$23 3 1 2 3 PMOS_VTG L=0.05U W=19.69U AS=2.22855P AD=2.22855P PS=25.565U
+ PD=25.565U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_13

* cell custom_sram_1r1w_32_256_freepdk45_pinv_12
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_12 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.26 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=2.16U AS=0.24705P AD=0.24705P PS=4.26U PD=4.26U
* device instance $9 r0 *1 0.2325,1.94 PMOS_VTG
M$9 3 1 2 3 PMOS_VTG L=0.05U W=6.48U AS=0.74115P AD=0.74115P PS=9.12U PD=9.12U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_12

* cell custom_sram_1r1w_32_256_freepdk45_pinv_11
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_11 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.245 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.72U AS=0.0846P AD=0.0846P PS=1.665U PD=1.665U
* device instance $4 r0 *1 0.2325,1.985 PMOS_VTG
M$4 3 1 2 3 PMOS_VTG L=0.05U W=2.16U AS=0.2538P AD=0.2538P PS=3.585U PD=3.585U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_11

* cell custom_sram_1r1w_32_256_freepdk45_pinv_10
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_10 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.26 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
* device instance $2 r0 *1 0.2325,1.94 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.81U AS=0.103275P AD=0.103275P PS=1.875U
+ PD=1.875U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_10

* cell custom_sram_1r1w_32_256_freepdk45_dff_buf_0
* pin Qb
* pin Q
* pin clk
* pin D
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_dff_buf_0 1 2 4 5 6 7
* net 1 Qb
* net 2 Q
* net 4 clk
* net 5 D
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 3.195,0
X$1 3 1 6 7 custom_sram_1r1w_32_256_freepdk45_pinv_5
* cell instance $2 r0 *1 3.8825,0
X$2 1 2 6 7 custom_sram_1r1w_32_256_freepdk45_pinv_6
* cell instance $5 r0 *1 0,0
X$5 3 5 4 6 7 dff
.ENDS custom_sram_1r1w_32_256_freepdk45_dff_buf_0

* cell custom_sram_1r1w_32_256_freepdk45_hierarchical_predecode2x4_0
* pin in_0
* pin in_1
* pin out_0
* pin out_1
* pin out_2
* pin out_3
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_hierarchical_predecode2x4_0 1 2 5 6 7
+ 8 9 10
* net 1 in_0
* net 2 in_1
* net 5 out_0
* net 6 out_1
* net 7 out_2
* net 8 out_3
* net 9 vdd
* net 10 gnd
* cell instance $1 r0 *1 0.56,0
X$1 1 3 9 10 custom_sram_1r1w_32_256_freepdk45_pinv_4
* cell instance $2 m0 *1 2.0875,4.94
X$2 6 1 4 9 10 custom_sram_1r1w_32_256_freepdk45_pand2
* cell instance $3 m0 *1 2.0875,9.88
X$3 8 1 2 9 10 custom_sram_1r1w_32_256_freepdk45_pand2
* cell instance $9 r0 *1 2.0875,4.94
X$9 7 3 2 9 10 custom_sram_1r1w_32_256_freepdk45_pand2
* cell instance $10 m0 *1 0.56,4.94
X$10 2 4 9 10 custom_sram_1r1w_32_256_freepdk45_pinv_4
* cell instance $16 r0 *1 2.0875,0
X$16 5 3 4 9 10 custom_sram_1r1w_32_256_freepdk45_pand2
.ENDS custom_sram_1r1w_32_256_freepdk45_hierarchical_predecode2x4_0

* cell custom_sram_1r1w_32_256_freepdk45_pinv_2
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_2 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.185 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.36U AS=0.0423P AD=0.0423P PS=1.185U PD=1.185U
* device instance $4 r0 *1 0.2325,1.19 PMOS_VTG
M$4 3 1 2 3 PMOS_VTG L=0.05U W=1.08U AS=0.1269P AD=0.1269P PS=2.145U PD=2.145U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_2

* cell custom_sram_1r1w_32_256_freepdk45_wordline_driver_array
* pin in_0
* pin wl_0
* pin in_1
* pin wl_1
* pin in_2
* pin wl_2
* pin in_3
* pin wl_3
* pin in_4
* pin wl_4
* pin in_5
* pin wl_5
* pin in_6
* pin wl_6
* pin in_7
* pin wl_7
* pin in_8
* pin wl_8
* pin in_9
* pin wl_9
* pin in_10
* pin wl_10
* pin in_11
* pin wl_11
* pin in_12
* pin wl_12
* pin in_13
* pin wl_13
* pin in_14
* pin wl_14
* pin in_15
* pin wl_15
* pin in_16
* pin wl_16
* pin in_17
* pin wl_17
* pin in_18
* pin wl_18
* pin in_19
* pin wl_19
* pin in_20
* pin wl_20
* pin in_21
* pin wl_21
* pin in_22
* pin wl_22
* pin in_23
* pin wl_23
* pin in_24
* pin wl_24
* pin in_25
* pin wl_25
* pin in_26
* pin wl_26
* pin in_27
* pin wl_27
* pin in_28
* pin wl_28
* pin in_29
* pin wl_29
* pin in_30
* pin wl_30
* pin in_31
* pin en
* pin wl_31
* pin in_32
* pin wl_32
* pin wl_33
* pin in_33
* pin in_34
* pin wl_34
* pin wl_35
* pin in_35
* pin in_36
* pin wl_36
* pin wl_37
* pin in_37
* pin in_38
* pin wl_38
* pin wl_39
* pin in_39
* pin in_40
* pin wl_40
* pin wl_41
* pin in_41
* pin in_42
* pin wl_42
* pin wl_43
* pin in_43
* pin in_44
* pin wl_44
* pin wl_45
* pin in_45
* pin in_46
* pin wl_46
* pin wl_47
* pin in_47
* pin in_48
* pin wl_48
* pin wl_49
* pin in_49
* pin in_50
* pin wl_50
* pin wl_51
* pin in_51
* pin in_52
* pin wl_52
* pin wl_53
* pin in_53
* pin in_54
* pin wl_54
* pin wl_55
* pin in_55
* pin in_56
* pin wl_56
* pin wl_57
* pin in_57
* pin in_58
* pin wl_58
* pin wl_59
* pin in_59
* pin in_60
* pin wl_60
* pin wl_61
* pin in_61
* pin in_62
* pin wl_62
* pin wl_63
* pin in_63
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_wordline_driver_array 1 2 3 4 5 6 7 8
+ 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34
+ 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86
+ 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108
+ 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127
+ 128 129 130 131
* net 1 in_0
* net 2 wl_0
* net 3 in_1
* net 4 wl_1
* net 5 in_2
* net 6 wl_2
* net 7 in_3
* net 8 wl_3
* net 9 in_4
* net 10 wl_4
* net 11 in_5
* net 12 wl_5
* net 13 in_6
* net 14 wl_6
* net 15 in_7
* net 16 wl_7
* net 17 in_8
* net 18 wl_8
* net 19 in_9
* net 20 wl_9
* net 21 in_10
* net 22 wl_10
* net 23 in_11
* net 24 wl_11
* net 25 in_12
* net 26 wl_12
* net 27 in_13
* net 28 wl_13
* net 29 in_14
* net 30 wl_14
* net 31 in_15
* net 32 wl_15
* net 33 in_16
* net 34 wl_16
* net 35 in_17
* net 36 wl_17
* net 37 in_18
* net 38 wl_18
* net 39 in_19
* net 40 wl_19
* net 41 in_20
* net 42 wl_20
* net 43 in_21
* net 44 wl_21
* net 45 in_22
* net 46 wl_22
* net 47 in_23
* net 48 wl_23
* net 49 in_24
* net 50 wl_24
* net 51 in_25
* net 52 wl_25
* net 53 in_26
* net 54 wl_26
* net 55 in_27
* net 56 wl_27
* net 57 in_28
* net 58 wl_28
* net 59 in_29
* net 60 wl_29
* net 61 in_30
* net 62 wl_30
* net 63 in_31
* net 64 en
* net 65 wl_31
* net 66 in_32
* net 67 wl_32
* net 68 wl_33
* net 69 in_33
* net 70 in_34
* net 71 wl_34
* net 72 wl_35
* net 73 in_35
* net 74 in_36
* net 75 wl_36
* net 76 wl_37
* net 77 in_37
* net 78 in_38
* net 79 wl_38
* net 80 wl_39
* net 81 in_39
* net 82 in_40
* net 83 wl_40
* net 84 wl_41
* net 85 in_41
* net 86 in_42
* net 87 wl_42
* net 88 wl_43
* net 89 in_43
* net 90 in_44
* net 91 wl_44
* net 92 wl_45
* net 93 in_45
* net 94 in_46
* net 95 wl_46
* net 96 wl_47
* net 97 in_47
* net 98 in_48
* net 99 wl_48
* net 100 wl_49
* net 101 in_49
* net 102 in_50
* net 103 wl_50
* net 104 wl_51
* net 105 in_51
* net 106 in_52
* net 107 wl_52
* net 108 wl_53
* net 109 in_53
* net 110 in_54
* net 111 wl_54
* net 112 wl_55
* net 113 in_55
* net 114 in_56
* net 115 wl_56
* net 116 wl_57
* net 117 in_57
* net 118 in_58
* net 119 wl_58
* net 120 wl_59
* net 121 in_59
* net 122 in_60
* net 123 wl_60
* net 124 wl_61
* net 125 in_61
* net 126 in_62
* net 127 wl_62
* net 128 wl_63
* net 129 in_63
* net 130 vdd
* net 131 gnd
* cell instance $1 r0 *1 0.56,0
X$1 2 1 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $2 m0 *1 0.56,2.99
X$2 4 3 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $3 r0 *1 0.56,2.99
X$3 6 5 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $4 m0 *1 0.56,5.98
X$4 8 7 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $5 r0 *1 0.56,5.98
X$5 10 9 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $6 m0 *1 0.56,8.97
X$6 12 11 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $7 r0 *1 0.56,8.97
X$7 14 13 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $8 m0 *1 0.56,11.96
X$8 16 15 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $9 r0 *1 0.56,11.96
X$9 18 17 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $10 m0 *1 0.56,14.95
X$10 20 19 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $11 r0 *1 0.56,14.95
X$11 22 21 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $12 m0 *1 0.56,17.94
X$12 24 23 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $13 r0 *1 0.56,17.94
X$13 26 25 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $14 m0 *1 0.56,20.93
X$14 28 27 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $15 r0 *1 0.56,20.93
X$15 30 29 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $16 m0 *1 0.56,23.92
X$16 32 31 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $17 r0 *1 0.56,23.92
X$17 34 33 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $18 m0 *1 0.56,26.91
X$18 36 35 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $19 r0 *1 0.56,26.91
X$19 38 37 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $20 m0 *1 0.56,29.9
X$20 40 39 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $21 r0 *1 0.56,29.9
X$21 42 41 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $22 m0 *1 0.56,32.89
X$22 44 43 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $23 r0 *1 0.56,32.89
X$23 46 45 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $24 m0 *1 0.56,35.88
X$24 48 47 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $25 r0 *1 0.56,35.88
X$25 50 49 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $26 m0 *1 0.56,38.87
X$26 52 51 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $27 r0 *1 0.56,38.87
X$27 54 53 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $28 m0 *1 0.56,41.86
X$28 56 55 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $29 r0 *1 0.56,41.86
X$29 58 57 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $30 m0 *1 0.56,44.85
X$30 60 59 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $31 r0 *1 0.56,44.85
X$31 62 61 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $32 m0 *1 0.56,47.84
X$32 65 63 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $34 m0 *1 0.56,80.73
X$34 108 109 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $36 r0 *1 0.56,80.73
X$36 111 110 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $38 m0 *1 0.56,95.68
X$38 128 129 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $42 r0 *1 0.56,77.74
X$42 107 106 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $49 m0 *1 0.56,83.72
X$49 112 113 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $52 r0 *1 0.56,71.76
X$52 99 98 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $54 m0 *1 0.56,74.75
X$54 100 101 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $56 r0 *1 0.56,74.75
X$56 103 102 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $59 m0 *1 0.56,77.74
X$59 104 105 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $65 r0 *1 0.56,86.71
X$65 119 118 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $67 m0 *1 0.56,86.71
X$67 116 117 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $69 r0 *1 0.56,92.69
X$69 127 126 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $71 m0 *1 0.56,92.69
X$71 124 125 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $73 r0 *1 0.56,89.7
X$73 123 122 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $75 m0 *1 0.56,89.7
X$75 120 121 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $77 r0 *1 0.56,83.72
X$77 115 114 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $84 m0 *1 0.56,59.8
X$84 80 81 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $93 r0 *1 0.56,56.81
X$93 79 78 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $95 m0 *1 0.56,56.81
X$95 76 77 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $97 r0 *1 0.56,53.82
X$97 75 74 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $99 m0 *1 0.56,53.82
X$99 72 73 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $101 r0 *1 0.56,50.83
X$101 71 70 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $103 m0 *1 0.56,50.83
X$103 68 69 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $105 r0 *1 0.56,47.84
X$105 67 66 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $114 m0 *1 0.56,71.76
X$114 96 97 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $116 r0 *1 0.56,68.77
X$116 95 94 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $118 r0 *1 0.56,65.78
X$118 91 90 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $120 m0 *1 0.56,65.78
X$120 88 89 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $122 r0 *1 0.56,62.79
X$122 87 86 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $124 m0 *1 0.56,62.79
X$124 84 85 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $126 r0 *1 0.56,59.8
X$126 83 82 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
* cell instance $128 m0 *1 0.56,68.77
X$128 92 93 64 130 131 custom_sram_1r1w_32_256_freepdk45_wordline_driver
.ENDS custom_sram_1r1w_32_256_freepdk45_wordline_driver_array

* cell custom_sram_1r1w_32_256_freepdk45_hierarchical_decoder
* pin decode_1
* pin decode_0
* pin addr_1
* pin addr_0
* pin decode_2
* pin decode_3
* pin decode_5
* pin decode_4
* pin decode_7
* pin decode_6
* pin addr_2
* pin addr_3
* pin addr_4
* pin addr_5
* pin decode_8
* pin decode_10
* pin decode_11
* pin decode_9
* pin decode_12
* pin decode_14
* pin decode_13
* pin decode_17
* pin decode_16
* pin decode_15
* pin decode_18
* pin decode_19
* pin decode_20
* pin decode_21
* pin decode_22
* pin decode_23
* pin decode_24
* pin decode_25
* pin decode_26
* pin decode_27
* pin decode_28
* pin decode_29
* pin decode_30
* pin decode_31
* pin decode_32
* pin decode_33
* pin decode_34
* pin decode_35
* pin decode_36
* pin decode_37
* pin decode_38
* pin decode_39
* pin decode_40
* pin decode_41
* pin decode_42
* pin decode_43
* pin decode_44
* pin decode_45
* pin decode_46
* pin decode_47
* pin decode_48
* pin decode_49
* pin decode_50
* pin decode_51
* pin decode_52
* pin decode_53
* pin decode_54
* pin decode_55
* pin decode_56
* pin decode_57
* pin decode_58
* pin decode_59
* pin decode_60
* pin decode_61
* pin decode_62
* pin decode_63
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_hierarchical_decoder 6 7 8 9 11 12 14
+ 15 17 18 19 20 21 22 24 25 26 27 29 32 33 34 35 36 37 38 39 40 41 42 43 44 45
+ 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71
+ 72 73 74 75 76 77 78 79 80 81 82 83 84
* net 6 decode_1
* net 7 decode_0
* net 8 addr_1
* net 9 addr_0
* net 11 decode_2
* net 12 decode_3
* net 14 decode_5
* net 15 decode_4
* net 17 decode_7
* net 18 decode_6
* net 19 addr_2
* net 20 addr_3
* net 21 addr_4
* net 22 addr_5
* net 24 decode_8
* net 25 decode_10
* net 26 decode_11
* net 27 decode_9
* net 29 decode_12
* net 32 decode_14
* net 33 decode_13
* net 34 decode_17
* net 35 decode_16
* net 36 decode_15
* net 37 decode_18
* net 38 decode_19
* net 39 decode_20
* net 40 decode_21
* net 41 decode_22
* net 42 decode_23
* net 43 decode_24
* net 44 decode_25
* net 45 decode_26
* net 46 decode_27
* net 47 decode_28
* net 48 decode_29
* net 49 decode_30
* net 50 decode_31
* net 51 decode_32
* net 52 decode_33
* net 53 decode_34
* net 54 decode_35
* net 55 decode_36
* net 56 decode_37
* net 57 decode_38
* net 58 decode_39
* net 59 decode_40
* net 60 decode_41
* net 61 decode_42
* net 62 decode_43
* net 63 decode_44
* net 64 decode_45
* net 65 decode_46
* net 66 decode_47
* net 67 decode_48
* net 68 decode_49
* net 69 decode_50
* net 70 decode_51
* net 71 decode_52
* net 72 decode_53
* net 73 decode_54
* net 74 decode_55
* net 75 decode_56
* net 76 decode_57
* net 77 decode_58
* net 78 decode_59
* net 79 decode_60
* net 80 decode_61
* net 81 decode_62
* net 82 decode_63
* net 83 vdd
* net 84 gnd
* cell instance $2 r0 *1 6.58,0
X$2 7 1 4 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $3 r0 *1 6.58,83.72
X$3 75 1 16 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $4 r0 *1 6.58,11.96
X$4 24 1 16 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $5 r0 *1 6.58,23.92
X$5 35 1 4 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $6 r0 *1 6.58,89.7
X$6 79 1 23 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $7 r0 *1 6.58,41.86
X$7 47 1 23 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $8 r0 *1 6.58,71.76
X$8 67 1 4 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $9 r0 *1 6.58,65.78
X$9 63 1 23 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $10 r0 *1 6.58,35.88
X$10 43 1 16 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $11 r0 *1 6.58,47.84
X$11 51 1 4 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $12 r0 *1 6.58,59.8
X$12 59 1 16 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $13 r0 *1 6.58,77.74
X$13 71 1 13 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $14 r0 *1 6.58,17.94
X$14 29 1 23 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $15 r0 *1 6.58,29.9
X$15 39 1 13 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $16 r0 *1 6.58,53.82
X$16 55 1 13 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $17 r0 *1 6.58,5.98
X$17 15 1 13 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $19 r0 *1 0.9425,0
X$19 9 8 1 2 3 10 83 84
+ custom_sram_1r1w_32_256_freepdk45_hierarchical_predecode2x4
* cell instance $37 m0 *1 6.58,2.99
X$37 6 2 4 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $38 m0 *1 6.58,8.97
X$38 14 2 13 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $39 m0 *1 6.58,68.77
X$39 64 2 23 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $40 m0 *1 6.58,26.91
X$40 34 2 4 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $41 m0 *1 6.58,74.75
X$41 68 2 4 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $42 m0 *1 6.58,32.89
X$42 40 2 13 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $43 m0 *1 6.58,80.73
X$43 72 2 13 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $44 m0 *1 6.58,14.95
X$44 27 2 16 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $45 m0 *1 6.58,20.93
X$45 33 2 23 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $46 m0 *1 6.58,44.85
X$46 48 2 23 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $47 m0 *1 6.58,50.83
X$47 52 2 4 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $48 m0 *1 6.58,38.87
X$48 44 2 16 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $49 m0 *1 6.58,56.81
X$49 56 2 13 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $50 m0 *1 6.58,62.79
X$50 60 2 16 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $51 m0 *1 6.58,92.69
X$51 80 2 23 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $52 m0 *1 6.58,86.71
X$52 76 2 16 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $72 r0 *1 6.58,2.99
X$72 11 3 4 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $73 r0 *1 6.58,26.91
X$73 37 3 4 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $74 r0 *1 6.58,14.95
X$74 25 3 16 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $75 r0 *1 6.58,20.93
X$75 32 3 23 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $76 r0 *1 6.58,38.87
X$76 45 3 16 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $77 r0 *1 6.58,44.85
X$77 49 3 23 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $78 r0 *1 6.58,86.71
X$78 77 3 16 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $79 r0 *1 6.58,62.79
X$79 61 3 16 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $80 r0 *1 6.58,68.77
X$80 65 3 23 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $81 r0 *1 6.58,74.75
X$81 69 3 4 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $82 r0 *1 6.58,56.81
X$82 57 3 13 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $83 r0 *1 6.58,80.73
X$83 73 3 13 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $84 r0 *1 6.58,92.69
X$84 81 3 23 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $85 r0 *1 6.58,32.89
X$85 41 3 13 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $86 r0 *1 6.58,50.83
X$86 53 3 4 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $87 r0 *1 6.58,8.97
X$87 18 3 13 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $107 m0 *1 6.58,5.98
X$107 12 10 4 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $108 m0 *1 6.58,29.9
X$108 38 10 4 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $109 m0 *1 6.58,77.74
X$109 70 10 4 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $110 m0 *1 6.58,53.82
X$110 54 10 4 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $113 r0 *1 0.9425,8.97
X$113 19 20 4 13 16 23 83 84
+ custom_sram_1r1w_32_256_freepdk45_hierarchical_predecode2x4
* cell instance $131 m0 *1 6.58,11.96
X$131 17 10 13 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $132 m0 *1 6.58,17.94
X$132 26 10 16 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $133 m0 *1 6.58,23.92
X$133 36 10 23 5 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $136 r0 *1 0.9425,17.94
X$136 21 22 5 28 30 31 83 84
+ custom_sram_1r1w_32_256_freepdk45_hierarchical_predecode2x4
* cell instance $158 m0 *1 6.58,59.8
X$158 58 10 13 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $159 m0 *1 6.58,83.72
X$159 74 10 13 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $160 m0 *1 6.58,71.76
X$160 66 10 23 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $161 m0 *1 6.58,65.78
X$161 62 10 16 30 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $162 m0 *1 6.58,41.86
X$162 46 10 16 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $163 m0 *1 6.58,35.88
X$163 42 10 13 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $164 m0 *1 6.58,95.68
X$164 82 10 23 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $165 m0 *1 6.58,47.84
X$165 50 10 23 28 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
* cell instance $166 m0 *1 6.58,89.7
X$166 78 10 16 31 83 84 custom_sram_1r1w_32_256_freepdk45_and3_dec
.ENDS custom_sram_1r1w_32_256_freepdk45_hierarchical_decoder

* cell custom_sram_1r1w_32_256_freepdk45_column_mux_array_0
* pin br_out_31
* pin br_out_30
* pin br_out_29
* pin br_out_28
* pin br_out_27
* pin br_out_26
* pin br_out_25
* pin br_out_24
* pin br_out_0
* pin br_out_23
* pin br_out_22
* pin br_out_21
* pin br_out_20
* pin br_out_19
* pin br_out_18
* pin br_out_17
* pin br_out_16
* pin br_out_15
* pin br_out_1
* pin br_out_14
* pin br_out_13
* pin br_out_12
* pin br_out_11
* pin br_out_10
* pin br_out_9
* pin br_out_8
* pin br_out_7
* pin br_out_6
* pin br_out_2
* pin br_out_5
* pin br_out_4
* pin br_out_3
* pin sel_0
* pin sel_1
* pin bl_out_31
* pin bl_out_0
* pin bl_out_30
* pin bl_out_29
* pin bl_out_28
* pin bl_out_27
* pin bl_out_1
* pin bl_out_26
* pin bl_out_25
* pin bl_out_24
* pin bl_out_2
* pin bl_out_23
* pin bl_out_22
* pin bl_out_21
* pin bl_out_20
* pin bl_out_3
* pin bl_out_19
* pin bl_out_18
* pin bl_out_17
* pin bl_out_4
* pin bl_out_16
* pin bl_out_15
* pin bl_out_14
* pin bl_out_13
* pin bl_out_5
* pin bl_out_12
* pin bl_out_11
* pin bl_out_10
* pin bl_out_6
* pin bl_out_9
* pin bl_out_8
* pin bl_out_7
* pin sel_2
* pin sel_3
* pin bl_0
* pin br_0
* pin bl_1
* pin br_1
* pin bl_2
* pin br_2
* pin bl_3
* pin br_3
* pin bl_4
* pin br_4
* pin bl_5
* pin br_5
* pin bl_6
* pin br_6
* pin bl_7
* pin br_7
* pin bl_8
* pin br_8
* pin bl_9
* pin br_9
* pin bl_10
* pin br_10
* pin bl_11
* pin br_11
* pin bl_12
* pin br_12
* pin bl_13
* pin br_13
* pin bl_14
* pin br_14
* pin bl_15
* pin br_15
* pin bl_16
* pin br_16
* pin bl_17
* pin br_17
* pin bl_18
* pin br_18
* pin bl_19
* pin br_19
* pin bl_20
* pin br_20
* pin bl_21
* pin br_21
* pin bl_22
* pin br_22
* pin bl_23
* pin br_23
* pin bl_24
* pin br_24
* pin bl_25
* pin br_25
* pin bl_26
* pin br_26
* pin bl_27
* pin br_27
* pin bl_28
* pin br_28
* pin bl_29
* pin br_29
* pin bl_30
* pin br_30
* pin bl_31
* pin br_31
* pin bl_32
* pin br_32
* pin bl_33
* pin br_33
* pin bl_34
* pin br_34
* pin bl_35
* pin br_35
* pin bl_36
* pin br_36
* pin bl_37
* pin br_37
* pin bl_38
* pin br_38
* pin bl_39
* pin br_39
* pin bl_40
* pin br_40
* pin bl_41
* pin br_41
* pin bl_42
* pin br_42
* pin bl_43
* pin br_43
* pin bl_44
* pin br_44
* pin bl_45
* pin br_45
* pin bl_46
* pin br_46
* pin bl_47
* pin br_47
* pin bl_48
* pin br_48
* pin bl_49
* pin br_49
* pin bl_50
* pin br_50
* pin bl_51
* pin br_51
* pin bl_52
* pin br_52
* pin bl_53
* pin br_53
* pin bl_54
* pin br_54
* pin bl_55
* pin br_55
* pin bl_56
* pin br_56
* pin bl_57
* pin br_57
* pin bl_58
* pin br_58
* pin bl_59
* pin br_59
* pin bl_60
* pin br_60
* pin bl_61
* pin br_61
* pin bl_62
* pin br_62
* pin bl_63
* pin br_63
* pin bl_64
* pin br_64
* pin bl_65
* pin br_65
* pin bl_66
* pin br_66
* pin bl_67
* pin br_67
* pin bl_68
* pin br_68
* pin bl_69
* pin br_69
* pin bl_70
* pin br_70
* pin bl_71
* pin br_71
* pin bl_72
* pin br_72
* pin bl_73
* pin br_73
* pin bl_74
* pin br_74
* pin bl_75
* pin br_75
* pin bl_76
* pin br_76
* pin bl_77
* pin br_77
* pin bl_78
* pin br_78
* pin bl_79
* pin br_79
* pin bl_80
* pin br_80
* pin bl_81
* pin br_81
* pin bl_82
* pin br_82
* pin bl_83
* pin br_83
* pin bl_84
* pin br_84
* pin bl_85
* pin br_85
* pin bl_86
* pin br_86
* pin bl_87
* pin br_87
* pin bl_88
* pin br_88
* pin bl_89
* pin br_89
* pin bl_90
* pin br_90
* pin bl_91
* pin br_91
* pin bl_92
* pin br_92
* pin bl_93
* pin br_93
* pin bl_94
* pin br_94
* pin bl_95
* pin br_95
* pin bl_96
* pin br_96
* pin bl_97
* pin br_97
* pin bl_98
* pin br_98
* pin bl_99
* pin br_99
* pin bl_100
* pin br_100
* pin bl_101
* pin br_101
* pin bl_102
* pin br_102
* pin bl_103
* pin br_103
* pin bl_104
* pin br_104
* pin bl_105
* pin br_105
* pin bl_106
* pin br_106
* pin bl_107
* pin br_107
* pin bl_108
* pin br_108
* pin bl_109
* pin br_109
* pin bl_110
* pin br_110
* pin bl_111
* pin br_111
* pin bl_112
* pin br_112
* pin bl_113
* pin br_113
* pin bl_114
* pin br_114
* pin bl_115
* pin br_115
* pin bl_116
* pin br_116
* pin bl_117
* pin br_117
* pin bl_118
* pin br_118
* pin bl_119
* pin br_119
* pin bl_120
* pin br_120
* pin bl_121
* pin br_121
* pin bl_122
* pin br_122
* pin bl_123
* pin br_123
* pin bl_124
* pin br_124
* pin bl_125
* pin br_125
* pin bl_126
* pin br_126
* pin bl_127
* pin br_127
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_column_mux_array_0 1 2 3 4 5 6 7 8 9
+ 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35
+ 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87
+ 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109
+ 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128
+ 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147
+ 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166
+ 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185
+ 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204
+ 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223
+ 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299
+ 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318
+ 319 320 321 322 323 324 325
* net 1 br_out_31
* net 2 br_out_30
* net 3 br_out_29
* net 4 br_out_28
* net 5 br_out_27
* net 6 br_out_26
* net 7 br_out_25
* net 8 br_out_24
* net 9 br_out_0
* net 10 br_out_23
* net 11 br_out_22
* net 12 br_out_21
* net 13 br_out_20
* net 14 br_out_19
* net 15 br_out_18
* net 16 br_out_17
* net 17 br_out_16
* net 18 br_out_15
* net 19 br_out_1
* net 20 br_out_14
* net 21 br_out_13
* net 22 br_out_12
* net 23 br_out_11
* net 24 br_out_10
* net 25 br_out_9
* net 26 br_out_8
* net 27 br_out_7
* net 28 br_out_6
* net 29 br_out_2
* net 30 br_out_5
* net 31 br_out_4
* net 32 br_out_3
* net 33 sel_0
* net 34 sel_1
* net 35 bl_out_31
* net 36 bl_out_0
* net 37 bl_out_30
* net 38 bl_out_29
* net 39 bl_out_28
* net 40 bl_out_27
* net 41 bl_out_1
* net 42 bl_out_26
* net 43 bl_out_25
* net 44 bl_out_24
* net 45 bl_out_2
* net 46 bl_out_23
* net 47 bl_out_22
* net 48 bl_out_21
* net 49 bl_out_20
* net 50 bl_out_3
* net 51 bl_out_19
* net 52 bl_out_18
* net 53 bl_out_17
* net 54 bl_out_4
* net 55 bl_out_16
* net 56 bl_out_15
* net 57 bl_out_14
* net 58 bl_out_13
* net 59 bl_out_5
* net 60 bl_out_12
* net 61 bl_out_11
* net 62 bl_out_10
* net 63 bl_out_6
* net 64 bl_out_9
* net 65 bl_out_8
* net 66 bl_out_7
* net 67 sel_2
* net 68 sel_3
* net 69 bl_0
* net 70 br_0
* net 71 bl_1
* net 72 br_1
* net 73 bl_2
* net 74 br_2
* net 75 bl_3
* net 76 br_3
* net 77 bl_4
* net 78 br_4
* net 79 bl_5
* net 80 br_5
* net 81 bl_6
* net 82 br_6
* net 83 bl_7
* net 84 br_7
* net 85 bl_8
* net 86 br_8
* net 87 bl_9
* net 88 br_9
* net 89 bl_10
* net 90 br_10
* net 91 bl_11
* net 92 br_11
* net 93 bl_12
* net 94 br_12
* net 95 bl_13
* net 96 br_13
* net 97 bl_14
* net 98 br_14
* net 99 bl_15
* net 100 br_15
* net 101 bl_16
* net 102 br_16
* net 103 bl_17
* net 104 br_17
* net 105 bl_18
* net 106 br_18
* net 107 bl_19
* net 108 br_19
* net 109 bl_20
* net 110 br_20
* net 111 bl_21
* net 112 br_21
* net 113 bl_22
* net 114 br_22
* net 115 bl_23
* net 116 br_23
* net 117 bl_24
* net 118 br_24
* net 119 bl_25
* net 120 br_25
* net 121 bl_26
* net 122 br_26
* net 123 bl_27
* net 124 br_27
* net 125 bl_28
* net 126 br_28
* net 127 bl_29
* net 128 br_29
* net 129 bl_30
* net 130 br_30
* net 131 bl_31
* net 132 br_31
* net 133 bl_32
* net 134 br_32
* net 135 bl_33
* net 136 br_33
* net 137 bl_34
* net 138 br_34
* net 139 bl_35
* net 140 br_35
* net 141 bl_36
* net 142 br_36
* net 143 bl_37
* net 144 br_37
* net 145 bl_38
* net 146 br_38
* net 147 bl_39
* net 148 br_39
* net 149 bl_40
* net 150 br_40
* net 151 bl_41
* net 152 br_41
* net 153 bl_42
* net 154 br_42
* net 155 bl_43
* net 156 br_43
* net 157 bl_44
* net 158 br_44
* net 159 bl_45
* net 160 br_45
* net 161 bl_46
* net 162 br_46
* net 163 bl_47
* net 164 br_47
* net 165 bl_48
* net 166 br_48
* net 167 bl_49
* net 168 br_49
* net 169 bl_50
* net 170 br_50
* net 171 bl_51
* net 172 br_51
* net 173 bl_52
* net 174 br_52
* net 175 bl_53
* net 176 br_53
* net 177 bl_54
* net 178 br_54
* net 179 bl_55
* net 180 br_55
* net 181 bl_56
* net 182 br_56
* net 183 bl_57
* net 184 br_57
* net 185 bl_58
* net 186 br_58
* net 187 bl_59
* net 188 br_59
* net 189 bl_60
* net 190 br_60
* net 191 bl_61
* net 192 br_61
* net 193 bl_62
* net 194 br_62
* net 195 bl_63
* net 196 br_63
* net 197 bl_64
* net 198 br_64
* net 199 bl_65
* net 200 br_65
* net 201 bl_66
* net 202 br_66
* net 203 bl_67
* net 204 br_67
* net 205 bl_68
* net 206 br_68
* net 207 bl_69
* net 208 br_69
* net 209 bl_70
* net 210 br_70
* net 211 bl_71
* net 212 br_71
* net 213 bl_72
* net 214 br_72
* net 215 bl_73
* net 216 br_73
* net 217 bl_74
* net 218 br_74
* net 219 bl_75
* net 220 br_75
* net 221 bl_76
* net 222 br_76
* net 223 bl_77
* net 224 br_77
* net 225 bl_78
* net 226 br_78
* net 227 bl_79
* net 228 br_79
* net 229 bl_80
* net 230 br_80
* net 231 bl_81
* net 232 br_81
* net 233 bl_82
* net 234 br_82
* net 235 bl_83
* net 236 br_83
* net 237 bl_84
* net 238 br_84
* net 239 bl_85
* net 240 br_85
* net 241 bl_86
* net 242 br_86
* net 243 bl_87
* net 244 br_87
* net 245 bl_88
* net 246 br_88
* net 247 bl_89
* net 248 br_89
* net 249 bl_90
* net 250 br_90
* net 251 bl_91
* net 252 br_91
* net 253 bl_92
* net 254 br_92
* net 255 bl_93
* net 256 br_93
* net 257 bl_94
* net 258 br_94
* net 259 bl_95
* net 260 br_95
* net 261 bl_96
* net 262 br_96
* net 263 bl_97
* net 264 br_97
* net 265 bl_98
* net 266 br_98
* net 267 bl_99
* net 268 br_99
* net 269 bl_100
* net 270 br_100
* net 271 bl_101
* net 272 br_101
* net 273 bl_102
* net 274 br_102
* net 275 bl_103
* net 276 br_103
* net 277 bl_104
* net 278 br_104
* net 279 bl_105
* net 280 br_105
* net 281 bl_106
* net 282 br_106
* net 283 bl_107
* net 284 br_107
* net 285 bl_108
* net 286 br_108
* net 287 bl_109
* net 288 br_109
* net 289 bl_110
* net 290 br_110
* net 291 bl_111
* net 292 br_111
* net 293 bl_112
* net 294 br_112
* net 295 bl_113
* net 296 br_113
* net 297 bl_114
* net 298 br_114
* net 299 bl_115
* net 300 br_115
* net 301 bl_116
* net 302 br_116
* net 303 bl_117
* net 304 br_117
* net 305 bl_118
* net 306 br_118
* net 307 bl_119
* net 308 br_119
* net 309 bl_120
* net 310 br_120
* net 311 bl_121
* net 312 br_121
* net 313 bl_122
* net 314 br_122
* net 315 bl_123
* net 316 br_123
* net 317 bl_124
* net 318 br_124
* net 319 bl_125
* net 320 br_125
* net 321 bl_126
* net 322 br_126
* net 323 bl_127
* net 324 br_127
* net 325 gnd
* cell instance $1 r0 *1 207.2325,0.91
X$1 33 317 1 35 318 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $2 r0 *1 208.4075,0.91
X$2 34 319 1 35 320 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $3 r0 *1 209.5825,0.91
X$3 67 321 1 35 322 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $4 r0 *1 210.7575,0.91
X$4 68 323 1 35 324 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $9 r0 *1 202.5325,0.91
X$9 33 309 2 37 310 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $10 r0 *1 203.7075,0.91
X$10 34 311 2 37 312 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $11 r0 *1 206.0575,0.91
X$11 68 315 2 37 316 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $12 r0 *1 204.8825,0.91
X$12 67 313 2 37 314 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $17 r0 *1 197.8325,0.91
X$17 33 301 3 38 302 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $18 r0 *1 199.0075,0.91
X$18 34 303 3 38 304 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $19 r0 *1 201.3575,0.91
X$19 68 307 3 38 308 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $20 r0 *1 200.1825,0.91
X$20 67 305 3 38 306 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $25 r0 *1 194.3075,0.91
X$25 34 295 4 39 296 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $26 r0 *1 195.4825,0.91
X$26 67 297 4 39 298 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $27 r0 *1 193.1325,0.91
X$27 33 293 4 39 294 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $28 r0 *1 196.6575,0.91
X$28 68 299 4 39 300 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $33 r0 *1 188.4325,0.91
X$33 33 285 5 40 286 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $34 r0 *1 189.6075,0.91
X$34 34 287 5 40 288 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $35 r0 *1 190.7825,0.91
X$35 67 289 5 40 290 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $36 r0 *1 191.9575,0.91
X$36 68 291 5 40 292 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $41 r0 *1 183.7325,0.91
X$41 33 277 6 42 278 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $42 r0 *1 184.9075,0.91
X$42 34 279 6 42 280 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $43 r0 *1 186.0825,0.91
X$43 67 281 6 42 282 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $44 r0 *1 187.2575,0.91
X$44 68 283 6 42 284 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $49 r0 *1 179.0325,0.91
X$49 33 269 7 43 270 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $50 r0 *1 180.2075,0.91
X$50 34 271 7 43 272 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $51 r0 *1 181.3825,0.91
X$51 67 273 7 43 274 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $52 r0 *1 182.5575,0.91
X$52 68 275 7 43 276 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $57 r0 *1 175.5075,0.91
X$57 34 263 8 44 264 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $58 r0 *1 176.6825,0.91
X$58 67 265 8 44 266 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $59 r0 *1 177.8575,0.91
X$59 68 267 8 44 268 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $60 r0 *1 174.3325,0.91
X$60 33 261 8 44 262 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $65 r0 *1 9.6175,0.91
X$65 33 69 9 36 70 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $66 r0 *1 13.1425,0.91
X$66 68 75 9 36 76 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $67 r0 *1 11.9675,0.91
X$67 67 73 9 36 74 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $68 r0 *1 10.7925,0.91
X$68 34 71 9 36 72 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $73 r0 *1 152.3275,0.91
X$73 33 253 10 46 254 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $74 r0 *1 153.5025,0.91
X$74 34 255 10 46 256 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $75 r0 *1 154.6775,0.91
X$75 67 257 10 46 258 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $76 r0 *1 155.8525,0.91
X$76 68 259 10 46 260 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $81 r0 *1 148.8025,0.91
X$81 34 247 11 47 248 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $82 r0 *1 149.9775,0.91
X$82 67 249 11 47 250 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $83 r0 *1 147.6275,0.91
X$83 33 245 11 47 246 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $84 r0 *1 151.1525,0.91
X$84 68 251 11 47 252 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $89 r0 *1 142.9275,0.91
X$89 33 237 12 48 238 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $90 r0 *1 144.1025,0.91
X$90 34 239 12 48 240 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $91 r0 *1 145.2775,0.91
X$91 67 241 12 48 242 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $92 r0 *1 146.4525,0.91
X$92 68 243 12 48 244 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $97 r0 *1 138.2275,0.91
X$97 33 229 13 49 230 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $98 r0 *1 140.5775,0.91
X$98 67 233 13 49 234 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $99 r0 *1 141.7525,0.91
X$99 68 235 13 49 236 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $100 r0 *1 139.4025,0.91
X$100 34 231 13 49 232 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $105 r0 *1 134.7025,0.91
X$105 34 223 14 51 224 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $106 r0 *1 135.8775,0.91
X$106 67 225 14 51 226 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $107 r0 *1 133.5275,0.91
X$107 33 221 14 51 222 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $108 r0 *1 137.0525,0.91
X$108 68 227 14 51 228 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $113 r0 *1 128.8275,0.91
X$113 33 213 15 52 214 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $114 r0 *1 130.0025,0.91
X$114 34 215 15 52 216 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $115 r0 *1 131.1775,0.91
X$115 67 217 15 52 218 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $116 r0 *1 132.3525,0.91
X$116 68 219 15 52 220 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $121 r0 *1 125.3025,0.91
X$121 34 207 16 53 208 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $122 r0 *1 126.4775,0.91
X$122 67 209 16 53 210 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $123 r0 *1 127.6525,0.91
X$123 68 211 16 53 212 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $124 r0 *1 124.1275,0.91
X$124 33 205 16 53 206 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $129 r0 *1 122.9525,0.91
X$129 68 203 17 55 204 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $130 r0 *1 121.7775,0.91
X$130 67 201 17 55 202 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $131 r0 *1 120.6025,0.91
X$131 34 199 17 55 200 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $132 r0 *1 119.4275,0.91
X$132 33 197 17 55 198 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $137 r0 *1 97.4225,0.91
X$137 33 189 18 56 190 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $138 r0 *1 98.5975,0.91
X$138 34 191 18 56 192 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $139 r0 *1 100.9475,0.91
X$139 68 195 18 56 196 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $140 r0 *1 99.7725,0.91
X$140 67 193 18 56 194 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $145 r0 *1 15.4925,0.91
X$145 34 79 19 41 80 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $146 r0 *1 14.3175,0.91
X$146 33 77 19 41 78 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $147 r0 *1 16.6675,0.91
X$147 67 81 19 41 82 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $148 r0 *1 17.8425,0.91
X$148 68 83 19 41 84 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $153 r0 *1 96.2475,0.91
X$153 68 187 20 57 188 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $154 r0 *1 95.0725,0.91
X$154 67 185 20 57 186 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $155 r0 *1 93.8975,0.91
X$155 34 183 20 57 184 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $156 r0 *1 92.7225,0.91
X$156 33 181 20 57 182 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $161 r0 *1 88.0225,0.91
X$161 33 173 21 58 174 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $162 r0 *1 91.5475,0.91
X$162 68 179 21 58 180 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $163 r0 *1 89.1975,0.91
X$163 34 175 21 58 176 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $164 r0 *1 90.3725,0.91
X$164 67 177 21 58 178 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $169 r0 *1 84.4975,0.91
X$169 34 167 22 60 168 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $170 r0 *1 83.3225,0.91
X$170 33 165 22 60 166 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $171 r0 *1 85.6725,0.91
X$171 67 169 22 60 170 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $172 r0 *1 86.8475,0.91
X$172 68 171 22 60 172 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $177 r0 *1 78.6225,0.91
X$177 33 157 23 61 158 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $178 r0 *1 79.7975,0.91
X$178 34 159 23 61 160 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $179 r0 *1 80.9725,0.91
X$179 67 161 23 61 162 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $180 r0 *1 82.1475,0.91
X$180 68 163 23 61 164 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $185 r0 *1 73.9225,0.91
X$185 33 149 24 62 150 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $186 r0 *1 75.0975,0.91
X$186 34 151 24 62 152 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $187 r0 *1 76.2725,0.91
X$187 67 153 24 62 154 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $188 r0 *1 77.4475,0.91
X$188 68 155 24 62 156 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $193 r0 *1 69.2225,0.91
X$193 33 141 25 64 142 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $194 r0 *1 70.3975,0.91
X$194 34 143 25 64 144 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $195 r0 *1 71.5725,0.91
X$195 67 145 25 64 146 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $196 r0 *1 72.7475,0.91
X$196 68 147 25 64 148 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $201 r0 *1 64.5225,0.91
X$201 33 133 26 65 134 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $202 r0 *1 66.8725,0.91
X$202 67 137 26 65 138 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $203 r0 *1 68.0475,0.91
X$203 68 139 26 65 140 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $204 r0 *1 65.6975,0.91
X$204 34 135 26 65 136 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $209 r0 *1 46.0425,0.91
X$209 68 131 27 66 132 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $210 r0 *1 44.8675,0.91
X$210 67 129 27 66 130 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $211 r0 *1 43.6925,0.91
X$211 34 127 27 66 128 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $212 r0 *1 42.5175,0.91
X$212 33 125 27 66 126 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $217 r0 *1 41.3425,0.91
X$217 68 123 28 63 124 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $218 r0 *1 40.1675,0.91
X$218 67 121 28 63 122 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $219 r0 *1 38.9925,0.91
X$219 34 119 28 63 120 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $220 r0 *1 37.8175,0.91
X$220 33 117 28 63 118 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $225 r0 *1 22.5425,0.91
X$225 68 91 29 45 92 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $226 r0 *1 21.3675,0.91
X$226 67 89 29 45 90 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $227 r0 *1 19.0175,0.91
X$227 33 85 29 45 86 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $228 r0 *1 20.1925,0.91
X$228 34 87 29 45 88 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $233 r0 *1 33.1175,0.91
X$233 33 109 30 59 110 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $234 r0 *1 36.6425,0.91
X$234 68 115 30 59 116 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $235 r0 *1 35.4675,0.91
X$235 67 113 30 59 114 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $236 r0 *1 34.2925,0.91
X$236 34 111 30 59 112 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $241 r0 *1 31.9425,0.91
X$241 68 107 31 54 108 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $242 r0 *1 30.7675,0.91
X$242 67 105 31 54 106 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $243 r0 *1 29.5925,0.91
X$243 34 103 31 54 104 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $244 r0 *1 28.4175,0.91
X$244 33 101 31 54 102 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $249 r0 *1 27.2425,0.91
X$249 68 99 32 50 100 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $250 r0 *1 24.8925,0.91
X$250 34 95 32 50 96 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $251 r0 *1 23.7175,0.91
X$251 33 93 32 50 94 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
* cell instance $252 r0 *1 26.0675,0.91
X$252 67 97 32 50 98 325 custom_sram_1r1w_32_256_freepdk45_column_mux_0
.ENDS custom_sram_1r1w_32_256_freepdk45_column_mux_array_0

* cell custom_sram_1r1w_32_256_freepdk45_sense_amp_array
* pin data_0
* pin data_1
* pin data_2
* pin data_3
* pin data_4
* pin data_5
* pin data_6
* pin data_7
* pin data_8
* pin data_9
* pin data_10
* pin data_11
* pin data_12
* pin data_13
* pin data_14
* pin data_15
* pin data_16
* pin data_17
* pin data_18
* pin data_19
* pin data_20
* pin data_21
* pin data_22
* pin data_23
* pin data_24
* pin data_25
* pin data_26
* pin data_27
* pin data_28
* pin data_29
* pin data_30
* pin data_31
* pin bl_0
* pin en
* pin br_0
* pin bl_1
* pin br_1
* pin bl_2
* pin br_2
* pin bl_3
* pin br_3
* pin bl_4
* pin br_4
* pin bl_5
* pin br_5
* pin bl_6
* pin br_6
* pin bl_7
* pin br_7
* pin bl_8
* pin br_8
* pin bl_9
* pin br_9
* pin bl_10
* pin br_10
* pin bl_11
* pin br_11
* pin bl_12
* pin br_12
* pin bl_13
* pin br_13
* pin bl_14
* pin br_14
* pin bl_15
* pin br_15
* pin bl_16
* pin br_16
* pin bl_17
* pin br_17
* pin bl_18
* pin br_18
* pin bl_19
* pin br_19
* pin bl_20
* pin br_20
* pin bl_21
* pin br_21
* pin bl_22
* pin br_22
* pin bl_23
* pin br_23
* pin bl_24
* pin br_24
* pin bl_25
* pin br_25
* pin bl_26
* pin br_26
* pin bl_27
* pin br_27
* pin bl_28
* pin br_28
* pin bl_29
* pin br_29
* pin bl_30
* pin br_30
* pin bl_31
* pin br_31
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_sense_amp_array 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36
+ 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99
* net 1 data_0
* net 2 data_1
* net 3 data_2
* net 4 data_3
* net 5 data_4
* net 6 data_5
* net 7 data_6
* net 8 data_7
* net 9 data_8
* net 10 data_9
* net 11 data_10
* net 12 data_11
* net 13 data_12
* net 14 data_13
* net 15 data_14
* net 16 data_15
* net 17 data_16
* net 18 data_17
* net 19 data_18
* net 20 data_19
* net 21 data_20
* net 22 data_21
* net 23 data_22
* net 24 data_23
* net 25 data_24
* net 26 data_25
* net 27 data_26
* net 28 data_27
* net 29 data_28
* net 30 data_29
* net 31 data_30
* net 32 data_31
* net 33 bl_0
* net 34 en
* net 35 br_0
* net 36 bl_1
* net 37 br_1
* net 38 bl_2
* net 39 br_2
* net 40 bl_3
* net 41 br_3
* net 42 bl_4
* net 43 br_4
* net 44 bl_5
* net 45 br_5
* net 46 bl_6
* net 47 br_6
* net 48 bl_7
* net 49 br_7
* net 50 bl_8
* net 51 br_8
* net 52 bl_9
* net 53 br_9
* net 54 bl_10
* net 55 br_10
* net 56 bl_11
* net 57 br_11
* net 58 bl_12
* net 59 br_12
* net 60 bl_13
* net 61 br_13
* net 62 bl_14
* net 63 br_14
* net 64 bl_15
* net 65 br_15
* net 66 bl_16
* net 67 br_16
* net 68 bl_17
* net 69 br_17
* net 70 bl_18
* net 71 br_18
* net 72 bl_19
* net 73 br_19
* net 74 bl_20
* net 75 br_20
* net 76 bl_21
* net 77 br_21
* net 78 bl_22
* net 79 br_22
* net 80 bl_23
* net 81 br_23
* net 82 bl_24
* net 83 br_24
* net 84 bl_25
* net 85 br_25
* net 86 bl_26
* net 87 br_26
* net 88 bl_27
* net 89 br_27
* net 90 bl_28
* net 91 br_28
* net 92 bl_29
* net 93 br_29
* net 94 bl_30
* net 95 br_30
* net 96 bl_31
* net 97 br_31
* net 98 vdd
* net 99 gnd
* cell instance $1 r0 *1 9.6175,0
X$1 35 1 33 34 98 99 sense_amp
* cell instance $2 r0 *1 14.3175,0
X$2 37 2 36 34 98 99 sense_amp
* cell instance $3 r0 *1 19.0175,0
X$3 39 3 38 34 98 99 sense_amp
* cell instance $4 r0 *1 23.7175,0
X$4 41 4 40 34 98 99 sense_amp
* cell instance $5 r0 *1 28.4175,0
X$5 43 5 42 34 98 99 sense_amp
* cell instance $6 r0 *1 33.1175,0
X$6 45 6 44 34 98 99 sense_amp
* cell instance $7 r0 *1 37.8175,0
X$7 47 7 46 34 98 99 sense_amp
* cell instance $8 r0 *1 42.5175,0
X$8 49 8 48 34 98 99 sense_amp
* cell instance $9 r0 *1 64.5225,0
X$9 51 9 50 34 98 99 sense_amp
* cell instance $10 r0 *1 69.2225,0
X$10 53 10 52 34 98 99 sense_amp
* cell instance $11 r0 *1 73.9225,0
X$11 55 11 54 34 98 99 sense_amp
* cell instance $12 r0 *1 78.6225,0
X$12 57 12 56 34 98 99 sense_amp
* cell instance $13 r0 *1 83.3225,0
X$13 59 13 58 34 98 99 sense_amp
* cell instance $14 r0 *1 88.0225,0
X$14 61 14 60 34 98 99 sense_amp
* cell instance $15 r0 *1 92.7225,0
X$15 63 15 62 34 98 99 sense_amp
* cell instance $16 r0 *1 97.4225,0
X$16 65 16 64 34 98 99 sense_amp
* cell instance $17 r0 *1 119.4275,0
X$17 67 17 66 34 98 99 sense_amp
* cell instance $18 r0 *1 124.1275,0
X$18 69 18 68 34 98 99 sense_amp
* cell instance $19 r0 *1 128.8275,0
X$19 71 19 70 34 98 99 sense_amp
* cell instance $20 r0 *1 133.5275,0
X$20 73 20 72 34 98 99 sense_amp
* cell instance $21 r0 *1 138.2275,0
X$21 75 21 74 34 98 99 sense_amp
* cell instance $22 r0 *1 142.9275,0
X$22 77 22 76 34 98 99 sense_amp
* cell instance $23 r0 *1 147.6275,0
X$23 79 23 78 34 98 99 sense_amp
* cell instance $24 r0 *1 152.3275,0
X$24 81 24 80 34 98 99 sense_amp
* cell instance $25 r0 *1 174.3325,0
X$25 83 25 82 34 98 99 sense_amp
* cell instance $26 r0 *1 179.0325,0
X$26 85 26 84 34 98 99 sense_amp
* cell instance $27 r0 *1 183.7325,0
X$27 87 27 86 34 98 99 sense_amp
* cell instance $28 r0 *1 188.4325,0
X$28 89 28 88 34 98 99 sense_amp
* cell instance $29 r0 *1 193.1325,0
X$29 91 29 90 34 98 99 sense_amp
* cell instance $30 r0 *1 197.8325,0
X$30 93 30 92 34 98 99 sense_amp
* cell instance $31 r0 *1 202.5325,0
X$31 95 31 94 34 98 99 sense_amp
* cell instance $32 r0 *1 207.2325,0
X$32 97 32 96 34 98 99 sense_amp
.ENDS custom_sram_1r1w_32_256_freepdk45_sense_amp_array

* cell custom_sram_1r1w_32_256_freepdk45_precharge_array_0
* pin en_bar
* pin bl_0
* pin br_0
* pin bl_1
* pin br_1
* pin bl_2
* pin br_2
* pin bl_3
* pin br_3
* pin bl_4
* pin br_4
* pin bl_5
* pin br_5
* pin bl_6
* pin br_6
* pin bl_7
* pin br_7
* pin bl_8
* pin br_8
* pin bl_9
* pin br_9
* pin bl_10
* pin br_10
* pin bl_11
* pin br_11
* pin bl_12
* pin br_12
* pin bl_13
* pin br_13
* pin bl_14
* pin br_14
* pin bl_15
* pin br_15
* pin bl_16
* pin br_16
* pin bl_17
* pin br_17
* pin bl_18
* pin br_18
* pin bl_19
* pin br_19
* pin bl_20
* pin br_20
* pin bl_21
* pin br_21
* pin bl_22
* pin br_22
* pin bl_23
* pin br_23
* pin bl_24
* pin br_24
* pin bl_25
* pin br_25
* pin bl_26
* pin br_26
* pin bl_27
* pin br_27
* pin bl_28
* pin br_28
* pin bl_29
* pin br_29
* pin bl_30
* pin br_30
* pin bl_31
* pin br_31
* pin bl_32
* pin br_32
* pin bl_33
* pin br_33
* pin bl_34
* pin br_34
* pin bl_35
* pin br_35
* pin bl_36
* pin br_36
* pin bl_37
* pin br_37
* pin bl_38
* pin br_38
* pin bl_39
* pin br_39
* pin bl_40
* pin br_40
* pin bl_41
* pin br_41
* pin bl_42
* pin br_42
* pin bl_43
* pin br_43
* pin bl_44
* pin br_44
* pin bl_45
* pin br_45
* pin bl_46
* pin br_46
* pin bl_47
* pin br_47
* pin bl_48
* pin br_48
* pin bl_49
* pin br_49
* pin bl_50
* pin br_50
* pin bl_51
* pin br_51
* pin bl_52
* pin br_52
* pin bl_53
* pin br_53
* pin bl_54
* pin br_54
* pin bl_55
* pin br_55
* pin bl_56
* pin br_56
* pin bl_57
* pin br_57
* pin bl_58
* pin br_58
* pin bl_59
* pin br_59
* pin bl_60
* pin br_60
* pin bl_61
* pin br_61
* pin bl_62
* pin br_62
* pin bl_63
* pin br_63
* pin bl_64
* pin br_64
* pin bl_65
* pin br_65
* pin bl_66
* pin br_66
* pin bl_67
* pin br_67
* pin bl_68
* pin br_68
* pin bl_69
* pin br_69
* pin bl_70
* pin br_70
* pin bl_71
* pin br_71
* pin bl_72
* pin br_72
* pin bl_73
* pin br_73
* pin bl_74
* pin br_74
* pin bl_75
* pin br_75
* pin bl_76
* pin br_76
* pin bl_77
* pin br_77
* pin bl_78
* pin br_78
* pin bl_79
* pin br_79
* pin bl_80
* pin br_80
* pin bl_81
* pin br_81
* pin bl_82
* pin br_82
* pin bl_83
* pin br_83
* pin bl_84
* pin br_84
* pin bl_85
* pin br_85
* pin bl_86
* pin br_86
* pin bl_87
* pin br_87
* pin bl_88
* pin br_88
* pin bl_89
* pin br_89
* pin bl_90
* pin br_90
* pin bl_91
* pin br_91
* pin bl_92
* pin br_92
* pin bl_93
* pin br_93
* pin bl_94
* pin br_94
* pin bl_95
* pin br_95
* pin bl_96
* pin br_96
* pin bl_97
* pin br_97
* pin bl_98
* pin br_98
* pin bl_99
* pin br_99
* pin bl_100
* pin br_100
* pin bl_101
* pin br_101
* pin bl_102
* pin br_102
* pin bl_103
* pin br_103
* pin bl_104
* pin br_104
* pin bl_105
* pin br_105
* pin bl_106
* pin br_106
* pin bl_107
* pin br_107
* pin bl_108
* pin br_108
* pin bl_109
* pin br_109
* pin bl_110
* pin br_110
* pin bl_111
* pin br_111
* pin bl_112
* pin br_112
* pin bl_113
* pin br_113
* pin bl_114
* pin br_114
* pin bl_115
* pin br_115
* pin bl_116
* pin br_116
* pin bl_117
* pin br_117
* pin bl_118
* pin br_118
* pin bl_119
* pin br_119
* pin bl_120
* pin br_120
* pin bl_121
* pin br_121
* pin bl_122
* pin br_122
* pin bl_123
* pin br_123
* pin bl_124
* pin br_124
* pin bl_125
* pin br_125
* pin bl_126
* pin br_126
* pin bl_127
* pin br_127
* pin bl_128
* pin br_128
* pin vdd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_precharge_array_0 1 2 3 4 5 6 7 8 9
+ 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35
+ 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87
+ 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109
+ 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128
+ 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147
+ 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166
+ 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185
+ 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204
+ 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223
+ 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
* net 1 en_bar
* net 2 bl_0
* net 3 br_0
* net 4 bl_1
* net 5 br_1
* net 6 bl_2
* net 7 br_2
* net 8 bl_3
* net 9 br_3
* net 10 bl_4
* net 11 br_4
* net 12 bl_5
* net 13 br_5
* net 14 bl_6
* net 15 br_6
* net 16 bl_7
* net 17 br_7
* net 18 bl_8
* net 19 br_8
* net 20 bl_9
* net 21 br_9
* net 22 bl_10
* net 23 br_10
* net 24 bl_11
* net 25 br_11
* net 26 bl_12
* net 27 br_12
* net 28 bl_13
* net 29 br_13
* net 30 bl_14
* net 31 br_14
* net 32 bl_15
* net 33 br_15
* net 34 bl_16
* net 35 br_16
* net 36 bl_17
* net 37 br_17
* net 38 bl_18
* net 39 br_18
* net 40 bl_19
* net 41 br_19
* net 42 bl_20
* net 43 br_20
* net 44 bl_21
* net 45 br_21
* net 46 bl_22
* net 47 br_22
* net 48 bl_23
* net 49 br_23
* net 50 bl_24
* net 51 br_24
* net 52 bl_25
* net 53 br_25
* net 54 bl_26
* net 55 br_26
* net 56 bl_27
* net 57 br_27
* net 58 bl_28
* net 59 br_28
* net 60 bl_29
* net 61 br_29
* net 62 bl_30
* net 63 br_30
* net 64 bl_31
* net 65 br_31
* net 66 bl_32
* net 67 br_32
* net 68 bl_33
* net 69 br_33
* net 70 bl_34
* net 71 br_34
* net 72 bl_35
* net 73 br_35
* net 74 bl_36
* net 75 br_36
* net 76 bl_37
* net 77 br_37
* net 78 bl_38
* net 79 br_38
* net 80 bl_39
* net 81 br_39
* net 82 bl_40
* net 83 br_40
* net 84 bl_41
* net 85 br_41
* net 86 bl_42
* net 87 br_42
* net 88 bl_43
* net 89 br_43
* net 90 bl_44
* net 91 br_44
* net 92 bl_45
* net 93 br_45
* net 94 bl_46
* net 95 br_46
* net 96 bl_47
* net 97 br_47
* net 98 bl_48
* net 99 br_48
* net 100 bl_49
* net 101 br_49
* net 102 bl_50
* net 103 br_50
* net 104 bl_51
* net 105 br_51
* net 106 bl_52
* net 107 br_52
* net 108 bl_53
* net 109 br_53
* net 110 bl_54
* net 111 br_54
* net 112 bl_55
* net 113 br_55
* net 114 bl_56
* net 115 br_56
* net 116 bl_57
* net 117 br_57
* net 118 bl_58
* net 119 br_58
* net 120 bl_59
* net 121 br_59
* net 122 bl_60
* net 123 br_60
* net 124 bl_61
* net 125 br_61
* net 126 bl_62
* net 127 br_62
* net 128 bl_63
* net 129 br_63
* net 130 bl_64
* net 131 br_64
* net 132 bl_65
* net 133 br_65
* net 134 bl_66
* net 135 br_66
* net 136 bl_67
* net 137 br_67
* net 138 bl_68
* net 139 br_68
* net 140 bl_69
* net 141 br_69
* net 142 bl_70
* net 143 br_70
* net 144 bl_71
* net 145 br_71
* net 146 bl_72
* net 147 br_72
* net 148 bl_73
* net 149 br_73
* net 150 bl_74
* net 151 br_74
* net 152 bl_75
* net 153 br_75
* net 154 bl_76
* net 155 br_76
* net 156 bl_77
* net 157 br_77
* net 158 bl_78
* net 159 br_78
* net 160 bl_79
* net 161 br_79
* net 162 bl_80
* net 163 br_80
* net 164 bl_81
* net 165 br_81
* net 166 bl_82
* net 167 br_82
* net 168 bl_83
* net 169 br_83
* net 170 bl_84
* net 171 br_84
* net 172 bl_85
* net 173 br_85
* net 174 bl_86
* net 175 br_86
* net 176 bl_87
* net 177 br_87
* net 178 bl_88
* net 179 br_88
* net 180 bl_89
* net 181 br_89
* net 182 bl_90
* net 183 br_90
* net 184 bl_91
* net 185 br_91
* net 186 bl_92
* net 187 br_92
* net 188 bl_93
* net 189 br_93
* net 190 bl_94
* net 191 br_94
* net 192 bl_95
* net 193 br_95
* net 194 bl_96
* net 195 br_96
* net 196 bl_97
* net 197 br_97
* net 198 bl_98
* net 199 br_98
* net 200 bl_99
* net 201 br_99
* net 202 bl_100
* net 203 br_100
* net 204 bl_101
* net 205 br_101
* net 206 bl_102
* net 207 br_102
* net 208 bl_103
* net 209 br_103
* net 210 bl_104
* net 211 br_104
* net 212 bl_105
* net 213 br_105
* net 214 bl_106
* net 215 br_106
* net 216 bl_107
* net 217 br_107
* net 218 bl_108
* net 219 br_108
* net 220 bl_109
* net 221 br_109
* net 222 bl_110
* net 223 br_110
* net 224 bl_111
* net 225 br_111
* net 226 bl_112
* net 227 br_112
* net 228 bl_113
* net 229 br_113
* net 230 bl_114
* net 231 br_114
* net 232 bl_115
* net 233 br_115
* net 234 bl_116
* net 235 br_116
* net 236 bl_117
* net 237 br_117
* net 238 bl_118
* net 239 br_118
* net 240 bl_119
* net 241 br_119
* net 242 bl_120
* net 243 br_120
* net 244 bl_121
* net 245 br_121
* net 246 bl_122
* net 247 br_122
* net 248 bl_123
* net 249 br_123
* net 250 bl_124
* net 251 br_124
* net 252 bl_125
* net 253 br_125
* net 254 bl_126
* net 255 br_126
* net 256 bl_127
* net 257 br_127
* net 258 bl_128
* net 259 br_128
* net 260 vdd
* cell instance $1 r0 *1 65.6975,0
X$1 1 68 69 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $2 r0 *1 64.5225,0
X$2 1 66 67 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $3 r0 *1 66.8725,0
X$3 1 70 71 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $4 r0 *1 68.0475,0
X$4 1 72 73 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $5 r0 *1 69.2225,0
X$5 1 74 75 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $6 r0 *1 70.3975,0
X$6 1 76 77 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $7 r0 *1 71.5725,0
X$7 1 78 79 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $8 r0 *1 72.7475,0
X$8 1 80 81 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $9 r0 *1 73.9225,0
X$9 1 82 83 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $10 r0 *1 75.0975,0
X$10 1 84 85 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $11 r0 *1 76.2725,0
X$11 1 86 87 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $12 r0 *1 77.4475,0
X$12 1 88 89 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $13 r0 *1 78.6225,0
X$13 1 90 91 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $14 r0 *1 79.7975,0
X$14 1 92 93 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $15 r0 *1 80.9725,0
X$15 1 94 95 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $16 r0 *1 82.1475,0
X$16 1 96 97 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $17 r0 *1 83.3225,0
X$17 1 98 99 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $18 r0 *1 84.4975,0
X$18 1 100 101 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $19 r0 *1 85.6725,0
X$19 1 102 103 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $20 r0 *1 86.8475,0
X$20 1 104 105 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $21 r0 *1 88.0225,0
X$21 1 106 107 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $22 r0 *1 89.1975,0
X$22 1 108 109 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $23 r0 *1 90.3725,0
X$23 1 110 111 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $24 r0 *1 91.5475,0
X$24 1 112 113 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $25 r0 *1 92.7225,0
X$25 1 114 115 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $26 r0 *1 93.8975,0
X$26 1 116 117 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $27 r0 *1 95.0725,0
X$27 1 118 119 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $28 r0 *1 96.2475,0
X$28 1 120 121 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $29 r0 *1 97.4225,0
X$29 1 122 123 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $30 r0 *1 98.5975,0
X$30 1 124 125 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $31 r0 *1 99.7725,0
X$31 1 126 127 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $32 r0 *1 100.9475,0
X$32 1 128 129 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $33 r0 *1 175.5075,0
X$33 1 196 197 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $34 r0 *1 174.3325,0
X$34 1 194 195 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $35 r0 *1 176.6825,0
X$35 1 198 199 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $36 r0 *1 177.8575,0
X$36 1 200 201 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $37 r0 *1 179.0325,0
X$37 1 202 203 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $38 r0 *1 180.2075,0
X$38 1 204 205 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $39 r0 *1 181.3825,0
X$39 1 206 207 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $40 r0 *1 182.5575,0
X$40 1 208 209 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $41 r0 *1 183.7325,0
X$41 1 210 211 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $42 r0 *1 184.9075,0
X$42 1 212 213 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $43 r0 *1 186.0825,0
X$43 1 214 215 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $44 r0 *1 187.2575,0
X$44 1 216 217 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $45 r0 *1 188.4325,0
X$45 1 218 219 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $46 r0 *1 189.6075,0
X$46 1 220 221 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $47 r0 *1 190.7825,0
X$47 1 222 223 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $48 r0 *1 191.9575,0
X$48 1 224 225 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $49 r0 *1 193.1325,0
X$49 1 226 227 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $50 r0 *1 194.3075,0
X$50 1 228 229 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $51 r0 *1 195.4825,0
X$51 1 230 231 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $52 r0 *1 196.6575,0
X$52 1 232 233 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $53 r0 *1 197.8325,0
X$53 1 234 235 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $54 r0 *1 199.0075,0
X$54 1 236 237 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $55 r0 *1 200.1825,0
X$55 1 238 239 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $56 r0 *1 201.3575,0
X$56 1 240 241 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $57 r0 *1 202.5325,0
X$57 1 242 243 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $58 r0 *1 203.7075,0
X$58 1 244 245 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $59 r0 *1 204.8825,0
X$59 1 246 247 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $60 r0 *1 206.0575,0
X$60 1 248 249 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $61 r0 *1 207.2325,0
X$61 1 250 251 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $62 r0 *1 208.4075,0
X$62 1 252 253 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $63 r0 *1 209.5825,0
X$63 1 254 255 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $64 r0 *1 210.7575,0
X$64 1 256 257 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $65 r0 *1 211.9325,0
X$65 1 258 259 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $66 r0 *1 120.6025,0
X$66 1 132 133 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $67 r0 *1 119.4275,0
X$67 1 130 131 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $68 r0 *1 121.7775,0
X$68 1 134 135 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $69 r0 *1 122.9525,0
X$69 1 136 137 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $70 r0 *1 124.1275,0
X$70 1 138 139 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $71 r0 *1 125.3025,0
X$71 1 140 141 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $72 r0 *1 126.4775,0
X$72 1 142 143 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $73 r0 *1 127.6525,0
X$73 1 144 145 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $74 r0 *1 128.8275,0
X$74 1 146 147 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $75 r0 *1 130.0025,0
X$75 1 148 149 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $76 r0 *1 131.1775,0
X$76 1 150 151 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $77 r0 *1 132.3525,0
X$77 1 152 153 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $78 r0 *1 133.5275,0
X$78 1 154 155 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $79 r0 *1 134.7025,0
X$79 1 156 157 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $80 r0 *1 135.8775,0
X$80 1 158 159 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $81 r0 *1 137.0525,0
X$81 1 160 161 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $82 r0 *1 138.2275,0
X$82 1 162 163 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $83 r0 *1 139.4025,0
X$83 1 164 165 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $84 r0 *1 140.5775,0
X$84 1 166 167 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $85 r0 *1 141.7525,0
X$85 1 168 169 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $86 r0 *1 142.9275,0
X$86 1 170 171 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $87 r0 *1 144.1025,0
X$87 1 172 173 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $88 r0 *1 145.2775,0
X$88 1 174 175 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $89 r0 *1 146.4525,0
X$89 1 176 177 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $90 r0 *1 147.6275,0
X$90 1 178 179 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $91 r0 *1 148.8025,0
X$91 1 180 181 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $92 r0 *1 149.9775,0
X$92 1 182 183 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $93 r0 *1 151.1525,0
X$93 1 184 185 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $94 r0 *1 152.3275,0
X$94 1 186 187 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $95 r0 *1 153.5025,0
X$95 1 188 189 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $96 r0 *1 154.6775,0
X$96 1 190 191 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $97 r0 *1 155.8525,0
X$97 1 192 193 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $98 r0 *1 9.6175,0
X$98 1 2 3 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $99 r0 *1 10.7925,0
X$99 1 4 5 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $100 r0 *1 11.9675,0
X$100 1 6 7 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $101 r0 *1 13.1425,0
X$101 1 8 9 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $102 r0 *1 14.3175,0
X$102 1 10 11 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $103 r0 *1 15.4925,0
X$103 1 12 13 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $104 r0 *1 16.6675,0
X$104 1 14 15 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $105 r0 *1 17.8425,0
X$105 1 16 17 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $106 r0 *1 19.0175,0
X$106 1 18 19 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $107 r0 *1 20.1925,0
X$107 1 20 21 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $108 r0 *1 21.3675,0
X$108 1 22 23 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $109 r0 *1 22.5425,0
X$109 1 24 25 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $110 r0 *1 23.7175,0
X$110 1 26 27 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $111 r0 *1 24.8925,0
X$111 1 28 29 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $112 r0 *1 26.0675,0
X$112 1 30 31 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $113 r0 *1 27.2425,0
X$113 1 32 33 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $114 r0 *1 28.4175,0
X$114 1 34 35 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $115 r0 *1 29.5925,0
X$115 1 36 37 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $116 r0 *1 30.7675,0
X$116 1 38 39 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $117 r0 *1 31.9425,0
X$117 1 40 41 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $118 r0 *1 33.1175,0
X$118 1 42 43 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $119 r0 *1 34.2925,0
X$119 1 44 45 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $120 r0 *1 35.4675,0
X$120 1 46 47 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $121 r0 *1 36.6425,0
X$121 1 48 49 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $122 r0 *1 37.8175,0
X$122 1 50 51 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $123 r0 *1 38.9925,0
X$123 1 52 53 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $124 r0 *1 40.1675,0
X$124 1 54 55 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $125 r0 *1 41.3425,0
X$125 1 56 57 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $126 r0 *1 42.5175,0
X$126 1 58 59 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $127 r0 *1 43.6925,0
X$127 1 60 61 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $128 r0 *1 44.8675,0
X$128 1 62 63 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
* cell instance $129 r0 *1 46.0425,0
X$129 1 64 65 260 custom_sram_1r1w_32_256_freepdk45_precharge_1
.ENDS custom_sram_1r1w_32_256_freepdk45_precharge_array_0

* cell custom_sram_1r1w_32_256_freepdk45_column_mux_array
* pin br_out_31
* pin br_out_30
* pin br_out_29
* pin br_out_28
* pin br_out_27
* pin br_out_26
* pin br_out_25
* pin br_out_24
* pin br_out_0
* pin br_out_23
* pin br_out_22
* pin br_out_21
* pin br_out_20
* pin br_out_19
* pin br_out_18
* pin br_out_17
* pin br_out_16
* pin br_out_15
* pin br_out_1
* pin br_out_14
* pin br_out_13
* pin br_out_12
* pin br_out_11
* pin br_out_10
* pin br_out_9
* pin br_out_8
* pin br_out_7
* pin br_out_6
* pin br_out_2
* pin br_out_5
* pin br_out_4
* pin br_out_3
* pin sel_0
* pin sel_1
* pin bl_out_31
* pin bl_out_0
* pin bl_out_30
* pin bl_out_29
* pin bl_out_28
* pin bl_out_27
* pin bl_out_1
* pin bl_out_26
* pin bl_out_25
* pin bl_out_24
* pin bl_out_2
* pin bl_out_23
* pin bl_out_22
* pin bl_out_21
* pin bl_out_20
* pin bl_out_3
* pin bl_out_19
* pin bl_out_18
* pin bl_out_17
* pin bl_out_4
* pin bl_out_16
* pin bl_out_15
* pin bl_out_14
* pin bl_out_13
* pin bl_out_5
* pin bl_out_12
* pin bl_out_11
* pin bl_out_10
* pin bl_out_6
* pin bl_out_9
* pin bl_out_8
* pin bl_out_7
* pin sel_2
* pin sel_3
* pin bl_0
* pin br_0
* pin bl_1
* pin br_1
* pin bl_2
* pin br_2
* pin bl_3
* pin br_3
* pin bl_4
* pin br_4
* pin bl_5
* pin br_5
* pin bl_6
* pin br_6
* pin bl_7
* pin br_7
* pin bl_8
* pin br_8
* pin bl_9
* pin br_9
* pin bl_10
* pin br_10
* pin bl_11
* pin br_11
* pin bl_12
* pin br_12
* pin bl_13
* pin br_13
* pin bl_14
* pin br_14
* pin bl_15
* pin br_15
* pin bl_16
* pin br_16
* pin bl_17
* pin br_17
* pin bl_18
* pin br_18
* pin bl_19
* pin br_19
* pin bl_20
* pin br_20
* pin bl_21
* pin br_21
* pin bl_22
* pin br_22
* pin bl_23
* pin br_23
* pin bl_24
* pin br_24
* pin bl_25
* pin br_25
* pin bl_26
* pin br_26
* pin bl_27
* pin br_27
* pin bl_28
* pin br_28
* pin bl_29
* pin br_29
* pin bl_30
* pin br_30
* pin bl_31
* pin br_31
* pin bl_32
* pin br_32
* pin bl_33
* pin br_33
* pin bl_34
* pin br_34
* pin bl_35
* pin br_35
* pin bl_36
* pin br_36
* pin bl_37
* pin br_37
* pin bl_38
* pin br_38
* pin bl_39
* pin br_39
* pin bl_40
* pin br_40
* pin bl_41
* pin br_41
* pin bl_42
* pin br_42
* pin bl_43
* pin br_43
* pin bl_44
* pin br_44
* pin bl_45
* pin br_45
* pin bl_46
* pin br_46
* pin bl_47
* pin br_47
* pin bl_48
* pin br_48
* pin bl_49
* pin br_49
* pin bl_50
* pin br_50
* pin bl_51
* pin br_51
* pin bl_52
* pin br_52
* pin bl_53
* pin br_53
* pin bl_54
* pin br_54
* pin bl_55
* pin br_55
* pin bl_56
* pin br_56
* pin bl_57
* pin br_57
* pin bl_58
* pin br_58
* pin bl_59
* pin br_59
* pin bl_60
* pin br_60
* pin bl_61
* pin br_61
* pin bl_62
* pin br_62
* pin bl_63
* pin br_63
* pin bl_64
* pin br_64
* pin bl_65
* pin br_65
* pin bl_66
* pin br_66
* pin bl_67
* pin br_67
* pin bl_68
* pin br_68
* pin bl_69
* pin br_69
* pin bl_70
* pin br_70
* pin bl_71
* pin br_71
* pin bl_72
* pin br_72
* pin bl_73
* pin br_73
* pin bl_74
* pin br_74
* pin bl_75
* pin br_75
* pin bl_76
* pin br_76
* pin bl_77
* pin br_77
* pin bl_78
* pin br_78
* pin bl_79
* pin br_79
* pin bl_80
* pin br_80
* pin bl_81
* pin br_81
* pin bl_82
* pin br_82
* pin bl_83
* pin br_83
* pin bl_84
* pin br_84
* pin bl_85
* pin br_85
* pin bl_86
* pin br_86
* pin bl_87
* pin br_87
* pin bl_88
* pin br_88
* pin bl_89
* pin br_89
* pin bl_90
* pin br_90
* pin bl_91
* pin br_91
* pin bl_92
* pin br_92
* pin bl_93
* pin br_93
* pin bl_94
* pin br_94
* pin bl_95
* pin br_95
* pin bl_96
* pin br_96
* pin bl_97
* pin br_97
* pin bl_98
* pin br_98
* pin bl_99
* pin br_99
* pin bl_100
* pin br_100
* pin bl_101
* pin br_101
* pin bl_102
* pin br_102
* pin bl_103
* pin br_103
* pin bl_104
* pin br_104
* pin bl_105
* pin br_105
* pin bl_106
* pin br_106
* pin bl_107
* pin br_107
* pin bl_108
* pin br_108
* pin bl_109
* pin br_109
* pin bl_110
* pin br_110
* pin bl_111
* pin br_111
* pin bl_112
* pin br_112
* pin bl_113
* pin br_113
* pin bl_114
* pin br_114
* pin bl_115
* pin br_115
* pin bl_116
* pin br_116
* pin bl_117
* pin br_117
* pin bl_118
* pin br_118
* pin bl_119
* pin br_119
* pin bl_120
* pin br_120
* pin bl_121
* pin br_121
* pin bl_122
* pin br_122
* pin bl_123
* pin br_123
* pin bl_124
* pin br_124
* pin bl_125
* pin br_125
* pin bl_126
* pin br_126
* pin bl_127
* pin br_127
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_column_mux_array 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36
+ 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129
+ 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148
+ 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167
+ 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186
+ 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205
+ 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224
+ 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243
+ 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262
+ 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319
+ 320 321 322 323 324 325
* net 1 br_out_31
* net 2 br_out_30
* net 3 br_out_29
* net 4 br_out_28
* net 5 br_out_27
* net 6 br_out_26
* net 7 br_out_25
* net 8 br_out_24
* net 9 br_out_0
* net 10 br_out_23
* net 11 br_out_22
* net 12 br_out_21
* net 13 br_out_20
* net 14 br_out_19
* net 15 br_out_18
* net 16 br_out_17
* net 17 br_out_16
* net 18 br_out_15
* net 19 br_out_1
* net 20 br_out_14
* net 21 br_out_13
* net 22 br_out_12
* net 23 br_out_11
* net 24 br_out_10
* net 25 br_out_9
* net 26 br_out_8
* net 27 br_out_7
* net 28 br_out_6
* net 29 br_out_2
* net 30 br_out_5
* net 31 br_out_4
* net 32 br_out_3
* net 33 sel_0
* net 34 sel_1
* net 35 bl_out_31
* net 36 bl_out_0
* net 37 bl_out_30
* net 38 bl_out_29
* net 39 bl_out_28
* net 40 bl_out_27
* net 41 bl_out_1
* net 42 bl_out_26
* net 43 bl_out_25
* net 44 bl_out_24
* net 45 bl_out_2
* net 46 bl_out_23
* net 47 bl_out_22
* net 48 bl_out_21
* net 49 bl_out_20
* net 50 bl_out_3
* net 51 bl_out_19
* net 52 bl_out_18
* net 53 bl_out_17
* net 54 bl_out_4
* net 55 bl_out_16
* net 56 bl_out_15
* net 57 bl_out_14
* net 58 bl_out_13
* net 59 bl_out_5
* net 60 bl_out_12
* net 61 bl_out_11
* net 62 bl_out_10
* net 63 bl_out_6
* net 64 bl_out_9
* net 65 bl_out_8
* net 66 bl_out_7
* net 67 sel_2
* net 68 sel_3
* net 69 bl_0
* net 70 br_0
* net 71 bl_1
* net 72 br_1
* net 73 bl_2
* net 74 br_2
* net 75 bl_3
* net 76 br_3
* net 77 bl_4
* net 78 br_4
* net 79 bl_5
* net 80 br_5
* net 81 bl_6
* net 82 br_6
* net 83 bl_7
* net 84 br_7
* net 85 bl_8
* net 86 br_8
* net 87 bl_9
* net 88 br_9
* net 89 bl_10
* net 90 br_10
* net 91 bl_11
* net 92 br_11
* net 93 bl_12
* net 94 br_12
* net 95 bl_13
* net 96 br_13
* net 97 bl_14
* net 98 br_14
* net 99 bl_15
* net 100 br_15
* net 101 bl_16
* net 102 br_16
* net 103 bl_17
* net 104 br_17
* net 105 bl_18
* net 106 br_18
* net 107 bl_19
* net 108 br_19
* net 109 bl_20
* net 110 br_20
* net 111 bl_21
* net 112 br_21
* net 113 bl_22
* net 114 br_22
* net 115 bl_23
* net 116 br_23
* net 117 bl_24
* net 118 br_24
* net 119 bl_25
* net 120 br_25
* net 121 bl_26
* net 122 br_26
* net 123 bl_27
* net 124 br_27
* net 125 bl_28
* net 126 br_28
* net 127 bl_29
* net 128 br_29
* net 129 bl_30
* net 130 br_30
* net 131 bl_31
* net 132 br_31
* net 133 bl_32
* net 134 br_32
* net 135 bl_33
* net 136 br_33
* net 137 bl_34
* net 138 br_34
* net 139 bl_35
* net 140 br_35
* net 141 bl_36
* net 142 br_36
* net 143 bl_37
* net 144 br_37
* net 145 bl_38
* net 146 br_38
* net 147 bl_39
* net 148 br_39
* net 149 bl_40
* net 150 br_40
* net 151 bl_41
* net 152 br_41
* net 153 bl_42
* net 154 br_42
* net 155 bl_43
* net 156 br_43
* net 157 bl_44
* net 158 br_44
* net 159 bl_45
* net 160 br_45
* net 161 bl_46
* net 162 br_46
* net 163 bl_47
* net 164 br_47
* net 165 bl_48
* net 166 br_48
* net 167 bl_49
* net 168 br_49
* net 169 bl_50
* net 170 br_50
* net 171 bl_51
* net 172 br_51
* net 173 bl_52
* net 174 br_52
* net 175 bl_53
* net 176 br_53
* net 177 bl_54
* net 178 br_54
* net 179 bl_55
* net 180 br_55
* net 181 bl_56
* net 182 br_56
* net 183 bl_57
* net 184 br_57
* net 185 bl_58
* net 186 br_58
* net 187 bl_59
* net 188 br_59
* net 189 bl_60
* net 190 br_60
* net 191 bl_61
* net 192 br_61
* net 193 bl_62
* net 194 br_62
* net 195 bl_63
* net 196 br_63
* net 197 bl_64
* net 198 br_64
* net 199 bl_65
* net 200 br_65
* net 201 bl_66
* net 202 br_66
* net 203 bl_67
* net 204 br_67
* net 205 bl_68
* net 206 br_68
* net 207 bl_69
* net 208 br_69
* net 209 bl_70
* net 210 br_70
* net 211 bl_71
* net 212 br_71
* net 213 bl_72
* net 214 br_72
* net 215 bl_73
* net 216 br_73
* net 217 bl_74
* net 218 br_74
* net 219 bl_75
* net 220 br_75
* net 221 bl_76
* net 222 br_76
* net 223 bl_77
* net 224 br_77
* net 225 bl_78
* net 226 br_78
* net 227 bl_79
* net 228 br_79
* net 229 bl_80
* net 230 br_80
* net 231 bl_81
* net 232 br_81
* net 233 bl_82
* net 234 br_82
* net 235 bl_83
* net 236 br_83
* net 237 bl_84
* net 238 br_84
* net 239 bl_85
* net 240 br_85
* net 241 bl_86
* net 242 br_86
* net 243 bl_87
* net 244 br_87
* net 245 bl_88
* net 246 br_88
* net 247 bl_89
* net 248 br_89
* net 249 bl_90
* net 250 br_90
* net 251 bl_91
* net 252 br_91
* net 253 bl_92
* net 254 br_92
* net 255 bl_93
* net 256 br_93
* net 257 bl_94
* net 258 br_94
* net 259 bl_95
* net 260 br_95
* net 261 bl_96
* net 262 br_96
* net 263 bl_97
* net 264 br_97
* net 265 bl_98
* net 266 br_98
* net 267 bl_99
* net 268 br_99
* net 269 bl_100
* net 270 br_100
* net 271 bl_101
* net 272 br_101
* net 273 bl_102
* net 274 br_102
* net 275 bl_103
* net 276 br_103
* net 277 bl_104
* net 278 br_104
* net 279 bl_105
* net 280 br_105
* net 281 bl_106
* net 282 br_106
* net 283 bl_107
* net 284 br_107
* net 285 bl_108
* net 286 br_108
* net 287 bl_109
* net 288 br_109
* net 289 bl_110
* net 290 br_110
* net 291 bl_111
* net 292 br_111
* net 293 bl_112
* net 294 br_112
* net 295 bl_113
* net 296 br_113
* net 297 bl_114
* net 298 br_114
* net 299 bl_115
* net 300 br_115
* net 301 bl_116
* net 302 br_116
* net 303 bl_117
* net 304 br_117
* net 305 bl_118
* net 306 br_118
* net 307 bl_119
* net 308 br_119
* net 309 bl_120
* net 310 br_120
* net 311 bl_121
* net 312 br_121
* net 313 bl_122
* net 314 br_122
* net 315 bl_123
* net 316 br_123
* net 317 bl_124
* net 318 br_124
* net 319 bl_125
* net 320 br_125
* net 321 bl_126
* net 322 br_126
* net 323 bl_127
* net 324 br_127
* net 325 gnd
* cell instance $1 r0 *1 210.7575,0.91
X$1 68 323 1 35 324 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $2 r0 *1 208.4075,0.91
X$2 34 319 1 35 320 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $3 r0 *1 207.2325,0.91
X$3 33 317 1 35 318 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $4 r0 *1 209.5825,0.91
X$4 67 321 1 35 322 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $9 r0 *1 202.5325,0.91
X$9 33 309 2 37 310 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $10 r0 *1 203.7075,0.91
X$10 34 311 2 37 312 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $11 r0 *1 204.8825,0.91
X$11 67 313 2 37 314 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $12 r0 *1 206.0575,0.91
X$12 68 315 2 37 316 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $17 r0 *1 200.1825,0.91
X$17 67 305 3 38 306 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $18 r0 *1 199.0075,0.91
X$18 34 303 3 38 304 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $19 r0 *1 201.3575,0.91
X$19 68 307 3 38 308 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $20 r0 *1 197.8325,0.91
X$20 33 301 3 38 302 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $25 r0 *1 194.3075,0.91
X$25 34 295 4 39 296 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $26 r0 *1 193.1325,0.91
X$26 33 293 4 39 294 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $27 r0 *1 195.4825,0.91
X$27 67 297 4 39 298 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $28 r0 *1 196.6575,0.91
X$28 68 299 4 39 300 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $33 r0 *1 191.9575,0.91
X$33 68 291 5 40 292 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $34 r0 *1 190.7825,0.91
X$34 67 289 5 40 290 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $35 r0 *1 188.4325,0.91
X$35 33 285 5 40 286 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $36 r0 *1 189.6075,0.91
X$36 34 287 5 40 288 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $41 r0 *1 186.0825,0.91
X$41 67 281 6 42 282 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $42 r0 *1 184.9075,0.91
X$42 34 279 6 42 280 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $43 r0 *1 187.2575,0.91
X$43 68 283 6 42 284 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $44 r0 *1 183.7325,0.91
X$44 33 277 6 42 278 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $49 r0 *1 182.5575,0.91
X$49 68 275 7 43 276 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $50 r0 *1 181.3825,0.91
X$50 67 273 7 43 274 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $51 r0 *1 180.2075,0.91
X$51 34 271 7 43 272 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $52 r0 *1 179.0325,0.91
X$52 33 269 7 43 270 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $57 r0 *1 177.8575,0.91
X$57 68 267 8 44 268 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $58 r0 *1 176.6825,0.91
X$58 67 265 8 44 266 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $59 r0 *1 175.5075,0.91
X$59 34 263 8 44 264 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $60 r0 *1 174.3325,0.91
X$60 33 261 8 44 262 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $65 r0 *1 9.6175,0.91
X$65 33 69 9 36 70 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $66 r0 *1 13.1425,0.91
X$66 68 75 9 36 76 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $67 r0 *1 11.9675,0.91
X$67 67 73 9 36 74 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $68 r0 *1 10.7925,0.91
X$68 34 71 9 36 72 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $73 r0 *1 154.6775,0.91
X$73 67 257 10 46 258 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $74 r0 *1 153.5025,0.91
X$74 34 255 10 46 256 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $75 r0 *1 152.3275,0.91
X$75 33 253 10 46 254 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $76 r0 *1 155.8525,0.91
X$76 68 259 10 46 260 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $81 r0 *1 149.9775,0.91
X$81 67 249 11 47 250 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $82 r0 *1 151.1525,0.91
X$82 68 251 11 47 252 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $83 r0 *1 148.8025,0.91
X$83 34 247 11 47 248 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $84 r0 *1 147.6275,0.91
X$84 33 245 11 47 246 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $89 r0 *1 146.4525,0.91
X$89 68 243 12 48 244 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $90 r0 *1 145.2775,0.91
X$90 67 241 12 48 242 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $91 r0 *1 144.1025,0.91
X$91 34 239 12 48 240 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $92 r0 *1 142.9275,0.91
X$92 33 237 12 48 238 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $97 r0 *1 141.7525,0.91
X$97 68 235 13 49 236 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $98 r0 *1 139.4025,0.91
X$98 34 231 13 49 232 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $99 r0 *1 138.2275,0.91
X$99 33 229 13 49 230 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $100 r0 *1 140.5775,0.91
X$100 67 233 13 49 234 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $105 r0 *1 137.0525,0.91
X$105 68 227 14 51 228 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $106 r0 *1 135.8775,0.91
X$106 67 225 14 51 226 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $107 r0 *1 133.5275,0.91
X$107 33 221 14 51 222 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $108 r0 *1 134.7025,0.91
X$108 34 223 14 51 224 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $113 r0 *1 132.3525,0.91
X$113 68 219 15 52 220 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $114 r0 *1 131.1775,0.91
X$114 67 217 15 52 218 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $115 r0 *1 130.0025,0.91
X$115 34 215 15 52 216 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $116 r0 *1 128.8275,0.91
X$116 33 213 15 52 214 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $121 r0 *1 124.1275,0.91
X$121 33 205 16 53 206 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $122 r0 *1 125.3025,0.91
X$122 34 207 16 53 208 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $123 r0 *1 126.4775,0.91
X$123 67 209 16 53 210 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $124 r0 *1 127.6525,0.91
X$124 68 211 16 53 212 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $129 r0 *1 122.9525,0.91
X$129 68 203 17 55 204 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $130 r0 *1 121.7775,0.91
X$130 67 201 17 55 202 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $131 r0 *1 120.6025,0.91
X$131 34 199 17 55 200 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $132 r0 *1 119.4275,0.91
X$132 33 197 17 55 198 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $137 r0 *1 100.9475,0.91
X$137 68 195 18 56 196 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $138 r0 *1 99.7725,0.91
X$138 67 193 18 56 194 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $139 r0 *1 98.5975,0.91
X$139 34 191 18 56 192 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $140 r0 *1 97.4225,0.91
X$140 33 189 18 56 190 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $145 r0 *1 15.4925,0.91
X$145 34 79 19 41 80 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $146 r0 *1 14.3175,0.91
X$146 33 77 19 41 78 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $147 r0 *1 17.8425,0.91
X$147 68 83 19 41 84 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $148 r0 *1 16.6675,0.91
X$148 67 81 19 41 82 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $153 r0 *1 96.2475,0.91
X$153 68 187 20 57 188 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $154 r0 *1 95.0725,0.91
X$154 67 185 20 57 186 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $155 r0 *1 93.8975,0.91
X$155 34 183 20 57 184 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $156 r0 *1 92.7225,0.91
X$156 33 181 20 57 182 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $161 r0 *1 91.5475,0.91
X$161 68 179 21 58 180 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $162 r0 *1 90.3725,0.91
X$162 67 177 21 58 178 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $163 r0 *1 89.1975,0.91
X$163 34 175 21 58 176 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $164 r0 *1 88.0225,0.91
X$164 33 173 21 58 174 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $169 r0 *1 84.4975,0.91
X$169 34 167 22 60 168 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $170 r0 *1 83.3225,0.91
X$170 33 165 22 60 166 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $171 r0 *1 85.6725,0.91
X$171 67 169 22 60 170 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $172 r0 *1 86.8475,0.91
X$172 68 171 22 60 172 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $177 r0 *1 78.6225,0.91
X$177 33 157 23 61 158 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $178 r0 *1 79.7975,0.91
X$178 34 159 23 61 160 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $179 r0 *1 80.9725,0.91
X$179 67 161 23 61 162 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $180 r0 *1 82.1475,0.91
X$180 68 163 23 61 164 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $185 r0 *1 75.0975,0.91
X$185 34 151 24 62 152 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $186 r0 *1 76.2725,0.91
X$186 67 153 24 62 154 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $187 r0 *1 73.9225,0.91
X$187 33 149 24 62 150 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $188 r0 *1 77.4475,0.91
X$188 68 155 24 62 156 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $193 r0 *1 71.5725,0.91
X$193 67 145 25 64 146 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $194 r0 *1 70.3975,0.91
X$194 34 143 25 64 144 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $195 r0 *1 69.2225,0.91
X$195 33 141 25 64 142 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $196 r0 *1 72.7475,0.91
X$196 68 147 25 64 148 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $201 r0 *1 68.0475,0.91
X$201 68 139 26 65 140 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $202 r0 *1 66.8725,0.91
X$202 67 137 26 65 138 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $203 r0 *1 64.5225,0.91
X$203 33 133 26 65 134 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $204 r0 *1 65.6975,0.91
X$204 34 135 26 65 136 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $209 r0 *1 46.0425,0.91
X$209 68 131 27 66 132 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $210 r0 *1 43.6925,0.91
X$210 34 127 27 66 128 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $211 r0 *1 44.8675,0.91
X$211 67 129 27 66 130 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $212 r0 *1 42.5175,0.91
X$212 33 125 27 66 126 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $217 r0 *1 40.1675,0.91
X$217 67 121 28 63 122 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $218 r0 *1 37.8175,0.91
X$218 33 117 28 63 118 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $219 r0 *1 38.9925,0.91
X$219 34 119 28 63 120 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $220 r0 *1 41.3425,0.91
X$220 68 123 28 63 124 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $225 r0 *1 20.1925,0.91
X$225 34 87 29 45 88 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $226 r0 *1 19.0175,0.91
X$226 33 85 29 45 86 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $227 r0 *1 22.5425,0.91
X$227 68 91 29 45 92 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $228 r0 *1 21.3675,0.91
X$228 67 89 29 45 90 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $233 r0 *1 35.4675,0.91
X$233 67 113 30 59 114 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $234 r0 *1 34.2925,0.91
X$234 34 111 30 59 112 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $235 r0 *1 33.1175,0.91
X$235 33 109 30 59 110 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $236 r0 *1 36.6425,0.91
X$236 68 115 30 59 116 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $241 r0 *1 28.4175,0.91
X$241 33 101 31 54 102 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $242 r0 *1 29.5925,0.91
X$242 34 103 31 54 104 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $243 r0 *1 30.7675,0.91
X$243 67 105 31 54 106 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $244 r0 *1 31.9425,0.91
X$244 68 107 31 54 108 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $249 r0 *1 23.7175,0.91
X$249 33 93 32 50 94 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $250 r0 *1 24.8925,0.91
X$250 34 95 32 50 96 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $251 r0 *1 26.0675,0.91
X$251 67 97 32 50 98 325 custom_sram_1r1w_32_256_freepdk45_column_mux
* cell instance $252 r0 *1 27.2425,0.91
X$252 68 99 32 50 100 325 custom_sram_1r1w_32_256_freepdk45_column_mux
.ENDS custom_sram_1r1w_32_256_freepdk45_column_mux_array

* cell custom_sram_1r1w_32_256_freepdk45_write_driver_array
* pin data_0
* pin data_1
* pin data_2
* pin data_3
* pin data_4
* pin data_5
* pin data_6
* pin data_7
* pin data_8
* pin data_9
* pin data_10
* pin data_11
* pin data_12
* pin data_13
* pin data_14
* pin data_15
* pin data_16
* pin data_17
* pin data_18
* pin data_19
* pin data_20
* pin data_21
* pin data_22
* pin data_23
* pin data_24
* pin data_25
* pin data_26
* pin data_27
* pin data_28
* pin data_29
* pin data_30
* pin data_31
* pin br_0
* pin br_1
* pin br_2
* pin br_3
* pin br_4
* pin br_5
* pin br_6
* pin br_7
* pin br_8
* pin br_9
* pin br_10
* pin br_11
* pin br_12
* pin br_13
* pin br_14
* pin br_15
* pin en
* pin br_16
* pin br_17
* pin br_18
* pin br_19
* pin br_20
* pin br_21
* pin br_22
* pin br_23
* pin br_24
* pin br_25
* pin br_26
* pin br_27
* pin br_28
* pin br_29
* pin br_30
* pin br_31
* pin bl_0
* pin bl_1
* pin bl_2
* pin bl_3
* pin bl_4
* pin bl_5
* pin bl_6
* pin bl_7
* pin bl_8
* pin bl_9
* pin bl_10
* pin bl_11
* pin bl_12
* pin bl_13
* pin bl_14
* pin bl_15
* pin bl_16
* pin bl_17
* pin bl_18
* pin bl_19
* pin bl_20
* pin bl_21
* pin bl_22
* pin bl_23
* pin bl_24
* pin bl_25
* pin bl_26
* pin bl_27
* pin bl_28
* pin bl_29
* pin bl_30
* pin bl_31
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_write_driver_array 1 2 3 4 5 6 7 8 9
+ 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35
+ 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87
+ 88 89 90 91 92 93 94 95 96 97 98 99
* net 1 data_0
* net 2 data_1
* net 3 data_2
* net 4 data_3
* net 5 data_4
* net 6 data_5
* net 7 data_6
* net 8 data_7
* net 9 data_8
* net 10 data_9
* net 11 data_10
* net 12 data_11
* net 13 data_12
* net 14 data_13
* net 15 data_14
* net 16 data_15
* net 17 data_16
* net 18 data_17
* net 19 data_18
* net 20 data_19
* net 21 data_20
* net 22 data_21
* net 23 data_22
* net 24 data_23
* net 25 data_24
* net 26 data_25
* net 27 data_26
* net 28 data_27
* net 29 data_28
* net 30 data_29
* net 31 data_30
* net 32 data_31
* net 33 br_0
* net 34 br_1
* net 35 br_2
* net 36 br_3
* net 37 br_4
* net 38 br_5
* net 39 br_6
* net 40 br_7
* net 41 br_8
* net 42 br_9
* net 43 br_10
* net 44 br_11
* net 45 br_12
* net 46 br_13
* net 47 br_14
* net 48 br_15
* net 49 en
* net 50 br_16
* net 51 br_17
* net 52 br_18
* net 53 br_19
* net 54 br_20
* net 55 br_21
* net 56 br_22
* net 57 br_23
* net 58 br_24
* net 59 br_25
* net 60 br_26
* net 61 br_27
* net 62 br_28
* net 63 br_29
* net 64 br_30
* net 65 br_31
* net 66 bl_0
* net 67 bl_1
* net 68 bl_2
* net 69 bl_3
* net 70 bl_4
* net 71 bl_5
* net 72 bl_6
* net 73 bl_7
* net 74 bl_8
* net 75 bl_9
* net 76 bl_10
* net 77 bl_11
* net 78 bl_12
* net 79 bl_13
* net 80 bl_14
* net 81 bl_15
* net 82 bl_16
* net 83 bl_17
* net 84 bl_18
* net 85 bl_19
* net 86 bl_20
* net 87 bl_21
* net 88 bl_22
* net 89 bl_23
* net 90 bl_24
* net 91 bl_25
* net 92 bl_26
* net 93 bl_27
* net 94 bl_28
* net 95 bl_29
* net 96 bl_30
* net 97 bl_31
* net 98 vdd
* net 99 gnd
* cell instance $1 r0 *1 9.6175,0
X$1 1 49 33 66 98 99 write_driver
* cell instance $2 r0 *1 14.3175,0
X$2 2 49 34 67 98 99 write_driver
* cell instance $3 r0 *1 19.0175,0
X$3 3 49 35 68 98 99 write_driver
* cell instance $4 r0 *1 23.7175,0
X$4 4 49 36 69 98 99 write_driver
* cell instance $5 r0 *1 28.4175,0
X$5 5 49 37 70 98 99 write_driver
* cell instance $6 r0 *1 33.1175,0
X$6 6 49 38 71 98 99 write_driver
* cell instance $7 r0 *1 37.8175,0
X$7 7 49 39 72 98 99 write_driver
* cell instance $8 r0 *1 42.5175,0
X$8 8 49 40 73 98 99 write_driver
* cell instance $9 r0 *1 64.5225,0
X$9 9 49 41 74 98 99 write_driver
* cell instance $10 r0 *1 69.2225,0
X$10 10 49 42 75 98 99 write_driver
* cell instance $11 r0 *1 73.9225,0
X$11 11 49 43 76 98 99 write_driver
* cell instance $12 r0 *1 78.6225,0
X$12 12 49 44 77 98 99 write_driver
* cell instance $13 r0 *1 83.3225,0
X$13 13 49 45 78 98 99 write_driver
* cell instance $14 r0 *1 88.0225,0
X$14 14 49 46 79 98 99 write_driver
* cell instance $15 r0 *1 92.7225,0
X$15 15 49 47 80 98 99 write_driver
* cell instance $16 r0 *1 97.4225,0
X$16 16 49 48 81 98 99 write_driver
* cell instance $17 r0 *1 119.4275,0
X$17 17 49 50 82 98 99 write_driver
* cell instance $18 r0 *1 124.1275,0
X$18 18 49 51 83 98 99 write_driver
* cell instance $19 r0 *1 128.8275,0
X$19 19 49 52 84 98 99 write_driver
* cell instance $20 r0 *1 133.5275,0
X$20 20 49 53 85 98 99 write_driver
* cell instance $21 r0 *1 138.2275,0
X$21 21 49 54 86 98 99 write_driver
* cell instance $22 r0 *1 142.9275,0
X$22 22 49 55 87 98 99 write_driver
* cell instance $23 r0 *1 147.6275,0
X$23 23 49 56 88 98 99 write_driver
* cell instance $24 r0 *1 152.3275,0
X$24 24 49 57 89 98 99 write_driver
* cell instance $25 r0 *1 174.3325,0
X$25 25 49 58 90 98 99 write_driver
* cell instance $26 r0 *1 179.0325,0
X$26 26 49 59 91 98 99 write_driver
* cell instance $27 r0 *1 183.7325,0
X$27 27 49 60 92 98 99 write_driver
* cell instance $28 r0 *1 188.4325,0
X$28 28 49 61 93 98 99 write_driver
* cell instance $29 r0 *1 193.1325,0
X$29 29 49 62 94 98 99 write_driver
* cell instance $30 r0 *1 197.8325,0
X$30 30 49 63 95 98 99 write_driver
* cell instance $31 r0 *1 202.5325,0
X$31 31 49 64 96 98 99 write_driver
* cell instance $32 r0 *1 207.2325,0
X$32 32 49 65 97 98 99 write_driver
.ENDS custom_sram_1r1w_32_256_freepdk45_write_driver_array

* cell custom_sram_1r1w_32_256_freepdk45_precharge_array
* pin en_bar
* pin bl_0
* pin br_0
* pin bl_1
* pin br_1
* pin bl_2
* pin br_2
* pin bl_3
* pin br_3
* pin bl_4
* pin br_4
* pin bl_5
* pin br_5
* pin bl_6
* pin br_6
* pin bl_7
* pin br_7
* pin bl_8
* pin br_8
* pin bl_9
* pin br_9
* pin bl_10
* pin br_10
* pin bl_11
* pin br_11
* pin bl_12
* pin br_12
* pin bl_13
* pin br_13
* pin bl_14
* pin br_14
* pin bl_15
* pin br_15
* pin bl_16
* pin br_16
* pin bl_17
* pin br_17
* pin bl_18
* pin br_18
* pin bl_19
* pin br_19
* pin bl_20
* pin br_20
* pin bl_21
* pin br_21
* pin bl_22
* pin br_22
* pin bl_23
* pin br_23
* pin bl_24
* pin br_24
* pin bl_25
* pin br_25
* pin bl_26
* pin br_26
* pin bl_27
* pin br_27
* pin bl_28
* pin br_28
* pin bl_29
* pin br_29
* pin bl_30
* pin br_30
* pin bl_31
* pin br_31
* pin bl_32
* pin br_32
* pin bl_33
* pin br_33
* pin bl_34
* pin br_34
* pin bl_35
* pin br_35
* pin bl_36
* pin br_36
* pin bl_37
* pin br_37
* pin bl_38
* pin br_38
* pin bl_39
* pin br_39
* pin bl_40
* pin br_40
* pin bl_41
* pin br_41
* pin bl_42
* pin br_42
* pin bl_43
* pin br_43
* pin bl_44
* pin br_44
* pin bl_45
* pin br_45
* pin bl_46
* pin br_46
* pin bl_47
* pin br_47
* pin bl_48
* pin br_48
* pin bl_49
* pin br_49
* pin bl_50
* pin br_50
* pin bl_51
* pin br_51
* pin bl_52
* pin br_52
* pin bl_53
* pin br_53
* pin bl_54
* pin br_54
* pin bl_55
* pin br_55
* pin bl_56
* pin br_56
* pin bl_57
* pin br_57
* pin bl_58
* pin br_58
* pin bl_59
* pin br_59
* pin bl_60
* pin br_60
* pin bl_61
* pin br_61
* pin bl_62
* pin br_62
* pin bl_63
* pin br_63
* pin bl_64
* pin br_64
* pin bl_65
* pin br_65
* pin bl_66
* pin br_66
* pin bl_67
* pin br_67
* pin bl_68
* pin br_68
* pin bl_69
* pin br_69
* pin bl_70
* pin br_70
* pin bl_71
* pin br_71
* pin bl_72
* pin br_72
* pin bl_73
* pin br_73
* pin bl_74
* pin br_74
* pin bl_75
* pin br_75
* pin bl_76
* pin br_76
* pin bl_77
* pin br_77
* pin bl_78
* pin br_78
* pin bl_79
* pin br_79
* pin bl_80
* pin br_80
* pin bl_81
* pin br_81
* pin bl_82
* pin br_82
* pin bl_83
* pin br_83
* pin bl_84
* pin br_84
* pin bl_85
* pin br_85
* pin bl_86
* pin br_86
* pin bl_87
* pin br_87
* pin bl_88
* pin br_88
* pin bl_89
* pin br_89
* pin bl_90
* pin br_90
* pin bl_91
* pin br_91
* pin bl_92
* pin br_92
* pin bl_93
* pin br_93
* pin bl_94
* pin br_94
* pin bl_95
* pin br_95
* pin bl_96
* pin br_96
* pin bl_97
* pin br_97
* pin bl_98
* pin br_98
* pin bl_99
* pin br_99
* pin bl_100
* pin br_100
* pin bl_101
* pin br_101
* pin bl_102
* pin br_102
* pin bl_103
* pin br_103
* pin bl_104
* pin br_104
* pin bl_105
* pin br_105
* pin bl_106
* pin br_106
* pin bl_107
* pin br_107
* pin bl_108
* pin br_108
* pin bl_109
* pin br_109
* pin bl_110
* pin br_110
* pin bl_111
* pin br_111
* pin bl_112
* pin br_112
* pin bl_113
* pin br_113
* pin bl_114
* pin br_114
* pin bl_115
* pin br_115
* pin bl_116
* pin br_116
* pin bl_117
* pin br_117
* pin bl_118
* pin br_118
* pin bl_119
* pin br_119
* pin bl_120
* pin br_120
* pin bl_121
* pin br_121
* pin bl_122
* pin br_122
* pin bl_123
* pin br_123
* pin bl_124
* pin br_124
* pin bl_125
* pin br_125
* pin bl_126
* pin br_126
* pin bl_127
* pin br_127
* pin bl_128
* pin br_128
* pin vdd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_precharge_array 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36
+ 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129
+ 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148
+ 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167
+ 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186
+ 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205
+ 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224
+ 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243
+ 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
* net 1 en_bar
* net 2 bl_0
* net 3 br_0
* net 4 bl_1
* net 5 br_1
* net 6 bl_2
* net 7 br_2
* net 8 bl_3
* net 9 br_3
* net 10 bl_4
* net 11 br_4
* net 12 bl_5
* net 13 br_5
* net 14 bl_6
* net 15 br_6
* net 16 bl_7
* net 17 br_7
* net 18 bl_8
* net 19 br_8
* net 20 bl_9
* net 21 br_9
* net 22 bl_10
* net 23 br_10
* net 24 bl_11
* net 25 br_11
* net 26 bl_12
* net 27 br_12
* net 28 bl_13
* net 29 br_13
* net 30 bl_14
* net 31 br_14
* net 32 bl_15
* net 33 br_15
* net 34 bl_16
* net 35 br_16
* net 36 bl_17
* net 37 br_17
* net 38 bl_18
* net 39 br_18
* net 40 bl_19
* net 41 br_19
* net 42 bl_20
* net 43 br_20
* net 44 bl_21
* net 45 br_21
* net 46 bl_22
* net 47 br_22
* net 48 bl_23
* net 49 br_23
* net 50 bl_24
* net 51 br_24
* net 52 bl_25
* net 53 br_25
* net 54 bl_26
* net 55 br_26
* net 56 bl_27
* net 57 br_27
* net 58 bl_28
* net 59 br_28
* net 60 bl_29
* net 61 br_29
* net 62 bl_30
* net 63 br_30
* net 64 bl_31
* net 65 br_31
* net 66 bl_32
* net 67 br_32
* net 68 bl_33
* net 69 br_33
* net 70 bl_34
* net 71 br_34
* net 72 bl_35
* net 73 br_35
* net 74 bl_36
* net 75 br_36
* net 76 bl_37
* net 77 br_37
* net 78 bl_38
* net 79 br_38
* net 80 bl_39
* net 81 br_39
* net 82 bl_40
* net 83 br_40
* net 84 bl_41
* net 85 br_41
* net 86 bl_42
* net 87 br_42
* net 88 bl_43
* net 89 br_43
* net 90 bl_44
* net 91 br_44
* net 92 bl_45
* net 93 br_45
* net 94 bl_46
* net 95 br_46
* net 96 bl_47
* net 97 br_47
* net 98 bl_48
* net 99 br_48
* net 100 bl_49
* net 101 br_49
* net 102 bl_50
* net 103 br_50
* net 104 bl_51
* net 105 br_51
* net 106 bl_52
* net 107 br_52
* net 108 bl_53
* net 109 br_53
* net 110 bl_54
* net 111 br_54
* net 112 bl_55
* net 113 br_55
* net 114 bl_56
* net 115 br_56
* net 116 bl_57
* net 117 br_57
* net 118 bl_58
* net 119 br_58
* net 120 bl_59
* net 121 br_59
* net 122 bl_60
* net 123 br_60
* net 124 bl_61
* net 125 br_61
* net 126 bl_62
* net 127 br_62
* net 128 bl_63
* net 129 br_63
* net 130 bl_64
* net 131 br_64
* net 132 bl_65
* net 133 br_65
* net 134 bl_66
* net 135 br_66
* net 136 bl_67
* net 137 br_67
* net 138 bl_68
* net 139 br_68
* net 140 bl_69
* net 141 br_69
* net 142 bl_70
* net 143 br_70
* net 144 bl_71
* net 145 br_71
* net 146 bl_72
* net 147 br_72
* net 148 bl_73
* net 149 br_73
* net 150 bl_74
* net 151 br_74
* net 152 bl_75
* net 153 br_75
* net 154 bl_76
* net 155 br_76
* net 156 bl_77
* net 157 br_77
* net 158 bl_78
* net 159 br_78
* net 160 bl_79
* net 161 br_79
* net 162 bl_80
* net 163 br_80
* net 164 bl_81
* net 165 br_81
* net 166 bl_82
* net 167 br_82
* net 168 bl_83
* net 169 br_83
* net 170 bl_84
* net 171 br_84
* net 172 bl_85
* net 173 br_85
* net 174 bl_86
* net 175 br_86
* net 176 bl_87
* net 177 br_87
* net 178 bl_88
* net 179 br_88
* net 180 bl_89
* net 181 br_89
* net 182 bl_90
* net 183 br_90
* net 184 bl_91
* net 185 br_91
* net 186 bl_92
* net 187 br_92
* net 188 bl_93
* net 189 br_93
* net 190 bl_94
* net 191 br_94
* net 192 bl_95
* net 193 br_95
* net 194 bl_96
* net 195 br_96
* net 196 bl_97
* net 197 br_97
* net 198 bl_98
* net 199 br_98
* net 200 bl_99
* net 201 br_99
* net 202 bl_100
* net 203 br_100
* net 204 bl_101
* net 205 br_101
* net 206 bl_102
* net 207 br_102
* net 208 bl_103
* net 209 br_103
* net 210 bl_104
* net 211 br_104
* net 212 bl_105
* net 213 br_105
* net 214 bl_106
* net 215 br_106
* net 216 bl_107
* net 217 br_107
* net 218 bl_108
* net 219 br_108
* net 220 bl_109
* net 221 br_109
* net 222 bl_110
* net 223 br_110
* net 224 bl_111
* net 225 br_111
* net 226 bl_112
* net 227 br_112
* net 228 bl_113
* net 229 br_113
* net 230 bl_114
* net 231 br_114
* net 232 bl_115
* net 233 br_115
* net 234 bl_116
* net 235 br_116
* net 236 bl_117
* net 237 br_117
* net 238 bl_118
* net 239 br_118
* net 240 bl_119
* net 241 br_119
* net 242 bl_120
* net 243 br_120
* net 244 bl_121
* net 245 br_121
* net 246 bl_122
* net 247 br_122
* net 248 bl_123
* net 249 br_123
* net 250 bl_124
* net 251 br_124
* net 252 bl_125
* net 253 br_125
* net 254 bl_126
* net 255 br_126
* net 256 bl_127
* net 257 br_127
* net 258 bl_128
* net 259 br_128
* net 260 vdd
* cell instance $1 r0 *1 8.4425,0
X$1 1 2 3 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $2 r0 *1 9.6175,0
X$2 1 4 5 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $3 r0 *1 10.7925,0
X$3 1 6 7 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $4 r0 *1 11.9675,0
X$4 1 8 9 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $5 r0 *1 13.1425,0
X$5 1 10 11 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $6 r0 *1 14.3175,0
X$6 1 12 13 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $7 r0 *1 15.4925,0
X$7 1 14 15 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $8 r0 *1 16.6675,0
X$8 1 16 17 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $9 r0 *1 17.8425,0
X$9 1 18 19 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $10 r0 *1 19.0175,0
X$10 1 20 21 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $11 r0 *1 20.1925,0
X$11 1 22 23 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $12 r0 *1 21.3675,0
X$12 1 24 25 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $13 r0 *1 22.5425,0
X$13 1 26 27 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $14 r0 *1 23.7175,0
X$14 1 28 29 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $15 r0 *1 24.8925,0
X$15 1 30 31 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $16 r0 *1 26.0675,0
X$16 1 32 33 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $17 r0 *1 27.2425,0
X$17 1 34 35 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $18 r0 *1 28.4175,0
X$18 1 36 37 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $19 r0 *1 29.5925,0
X$19 1 38 39 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $20 r0 *1 30.7675,0
X$20 1 40 41 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $21 r0 *1 31.9425,0
X$21 1 42 43 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $22 r0 *1 33.1175,0
X$22 1 44 45 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $23 r0 *1 34.2925,0
X$23 1 46 47 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $24 r0 *1 35.4675,0
X$24 1 48 49 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $25 r0 *1 36.6425,0
X$25 1 50 51 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $26 r0 *1 37.8175,0
X$26 1 52 53 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $27 r0 *1 38.9925,0
X$27 1 54 55 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $28 r0 *1 40.1675,0
X$28 1 56 57 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $29 r0 *1 41.3425,0
X$29 1 58 59 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $30 r0 *1 42.5175,0
X$30 1 60 61 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $31 r0 *1 43.6925,0
X$31 1 62 63 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $32 r0 *1 44.8675,0
X$32 1 64 65 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $33 r0 *1 46.0425,0
X$33 1 66 67 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $34 r0 *1 65.6975,0
X$34 1 70 71 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $35 r0 *1 64.5225,0
X$35 1 68 69 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $36 r0 *1 66.8725,0
X$36 1 72 73 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $37 r0 *1 68.0475,0
X$37 1 74 75 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $38 r0 *1 69.2225,0
X$38 1 76 77 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $39 r0 *1 70.3975,0
X$39 1 78 79 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $40 r0 *1 71.5725,0
X$40 1 80 81 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $41 r0 *1 72.7475,0
X$41 1 82 83 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $42 r0 *1 73.9225,0
X$42 1 84 85 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $43 r0 *1 75.0975,0
X$43 1 86 87 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $44 r0 *1 76.2725,0
X$44 1 88 89 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $45 r0 *1 77.4475,0
X$45 1 90 91 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $46 r0 *1 78.6225,0
X$46 1 92 93 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $47 r0 *1 79.7975,0
X$47 1 94 95 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $48 r0 *1 80.9725,0
X$48 1 96 97 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $49 r0 *1 82.1475,0
X$49 1 98 99 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $50 r0 *1 83.3225,0
X$50 1 100 101 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $51 r0 *1 84.4975,0
X$51 1 102 103 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $52 r0 *1 85.6725,0
X$52 1 104 105 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $53 r0 *1 86.8475,0
X$53 1 106 107 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $54 r0 *1 88.0225,0
X$54 1 108 109 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $55 r0 *1 89.1975,0
X$55 1 110 111 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $56 r0 *1 90.3725,0
X$56 1 112 113 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $57 r0 *1 91.5475,0
X$57 1 114 115 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $58 r0 *1 92.7225,0
X$58 1 116 117 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $59 r0 *1 93.8975,0
X$59 1 118 119 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $60 r0 *1 95.0725,0
X$60 1 120 121 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $61 r0 *1 96.2475,0
X$61 1 122 123 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $62 r0 *1 97.4225,0
X$62 1 124 125 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $63 r0 *1 98.5975,0
X$63 1 126 127 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $64 r0 *1 99.7725,0
X$64 1 128 129 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $65 r0 *1 100.9475,0
X$65 1 130 131 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $66 r0 *1 120.6025,0
X$66 1 134 135 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $67 r0 *1 119.4275,0
X$67 1 132 133 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $68 r0 *1 121.7775,0
X$68 1 136 137 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $69 r0 *1 122.9525,0
X$69 1 138 139 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $70 r0 *1 124.1275,0
X$70 1 140 141 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $71 r0 *1 125.3025,0
X$71 1 142 143 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $72 r0 *1 126.4775,0
X$72 1 144 145 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $73 r0 *1 127.6525,0
X$73 1 146 147 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $74 r0 *1 128.8275,0
X$74 1 148 149 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $75 r0 *1 130.0025,0
X$75 1 150 151 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $76 r0 *1 131.1775,0
X$76 1 152 153 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $77 r0 *1 132.3525,0
X$77 1 154 155 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $78 r0 *1 133.5275,0
X$78 1 156 157 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $79 r0 *1 134.7025,0
X$79 1 158 159 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $80 r0 *1 135.8775,0
X$80 1 160 161 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $81 r0 *1 137.0525,0
X$81 1 162 163 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $82 r0 *1 138.2275,0
X$82 1 164 165 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $83 r0 *1 139.4025,0
X$83 1 166 167 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $84 r0 *1 140.5775,0
X$84 1 168 169 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $85 r0 *1 141.7525,0
X$85 1 170 171 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $86 r0 *1 142.9275,0
X$86 1 172 173 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $87 r0 *1 144.1025,0
X$87 1 174 175 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $88 r0 *1 145.2775,0
X$88 1 176 177 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $89 r0 *1 146.4525,0
X$89 1 178 179 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $90 r0 *1 147.6275,0
X$90 1 180 181 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $91 r0 *1 148.8025,0
X$91 1 182 183 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $92 r0 *1 149.9775,0
X$92 1 184 185 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $93 r0 *1 151.1525,0
X$93 1 186 187 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $94 r0 *1 152.3275,0
X$94 1 188 189 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $95 r0 *1 153.5025,0
X$95 1 190 191 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $96 r0 *1 154.6775,0
X$96 1 192 193 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $97 r0 *1 155.8525,0
X$97 1 194 195 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $98 r0 *1 175.5075,0
X$98 1 198 199 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $99 r0 *1 174.3325,0
X$99 1 196 197 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $100 r0 *1 176.6825,0
X$100 1 200 201 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $101 r0 *1 177.8575,0
X$101 1 202 203 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $102 r0 *1 179.0325,0
X$102 1 204 205 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $103 r0 *1 180.2075,0
X$103 1 206 207 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $104 r0 *1 181.3825,0
X$104 1 208 209 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $105 r0 *1 182.5575,0
X$105 1 210 211 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $106 r0 *1 183.7325,0
X$106 1 212 213 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $107 r0 *1 184.9075,0
X$107 1 214 215 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $108 r0 *1 186.0825,0
X$108 1 216 217 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $109 r0 *1 187.2575,0
X$109 1 218 219 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $110 r0 *1 188.4325,0
X$110 1 220 221 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $111 r0 *1 189.6075,0
X$111 1 222 223 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $112 r0 *1 190.7825,0
X$112 1 224 225 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $113 r0 *1 191.9575,0
X$113 1 226 227 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $114 r0 *1 193.1325,0
X$114 1 228 229 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $115 r0 *1 194.3075,0
X$115 1 230 231 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $116 r0 *1 195.4825,0
X$116 1 232 233 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $117 r0 *1 196.6575,0
X$117 1 234 235 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $118 r0 *1 197.8325,0
X$118 1 236 237 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $119 r0 *1 199.0075,0
X$119 1 238 239 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $120 r0 *1 200.1825,0
X$120 1 240 241 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $121 r0 *1 201.3575,0
X$121 1 242 243 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $122 r0 *1 202.5325,0
X$122 1 244 245 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $123 r0 *1 203.7075,0
X$123 1 246 247 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $124 r0 *1 204.8825,0
X$124 1 248 249 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $125 r0 *1 206.0575,0
X$125 1 250 251 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $126 r0 *1 207.2325,0
X$126 1 252 253 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $127 r0 *1 208.4075,0
X$127 1 254 255 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $128 r0 *1 209.5825,0
X$128 1 256 257 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
* cell instance $129 r0 *1 210.7575,0
X$129 1 258 259 260 custom_sram_1r1w_32_256_freepdk45_precharge_0
.ENDS custom_sram_1r1w_32_256_freepdk45_precharge_array

* cell custom_sram_1r1w_32_256_freepdk45_local_bitcell_array_1
* pin wl_0_3
* pin wl_0_4
* pin rbl_wl_0_0
* pin wl_0_1
* pin wl_0_0
* pin wl_0_6
* pin wl_0_2
* pin wl_0_5
* pin wl_1_1
* pin wl_1_0
* pin wl_1_6
* pin wl_1_2
* pin wl_1_4
* pin wl_1_3
* pin wl_1_5
* pin wl_0_9
* pin wl_0_10
* pin wl_0_8
* pin wl_0_11
* pin wl_0_12
* pin wl_0_7
* pin wl_0_13
* pin wl_0_14
* pin wl_1_7
* pin wl_1_13
* pin wl_1_8
* pin wl_1_9
* pin wl_1_10
* pin wl_1_11
* pin wl_1_12
* pin wl_0_20
* pin wl_0_17
* pin wl_0_16
* pin wl_0_18
* pin wl_0_19
* pin wl_0_15
* pin wl_0_21
* pin wl_1_15
* pin wl_1_14
* pin wl_1_21
* pin wl_1_18
* pin wl_1_19
* pin wl_1_17
* pin wl_1_16
* pin wl_1_20
* pin wl_0_27
* pin wl_0_24
* pin wl_0_28
* pin wl_0_23
* pin wl_0_29
* pin wl_0_22
* pin wl_0_26
* pin wl_0_25
* pin wl_1_24
* pin wl_1_22
* pin wl_1_27
* pin wl_1_28
* pin wl_1_25
* pin wl_1_26
* pin wl_1_23
* pin wl_0_30
* pin wl_0_31
* pin bl_0_0
* pin bl_1_0
* pin br_1_0
* pin br_0_0
* pin bl_0_1
* pin bl_1_1
* pin br_1_1
* pin br_0_1
* pin bl_0_2
* pin bl_1_2
* pin br_1_2
* pin br_0_2
* pin bl_0_3
* pin bl_1_3
* pin br_1_3
* pin br_0_3
* pin bl_0_4
* pin bl_1_4
* pin br_1_4
* pin br_0_4
* pin bl_0_5
* pin bl_1_5
* pin br_1_5
* pin br_0_5
* pin bl_0_6
* pin bl_1_6
* pin br_1_6
* pin br_0_6
* pin bl_0_7
* pin bl_1_7
* pin br_1_7
* pin br_0_7
* pin bl_0_8
* pin bl_1_8
* pin br_1_8
* pin br_0_8
* pin bl_0_9
* pin bl_1_9
* pin br_1_9
* pin br_0_9
* pin bl_0_10
* pin bl_1_10
* pin br_1_10
* pin br_0_10
* pin bl_0_11
* pin bl_1_11
* pin br_1_11
* pin br_0_11
* pin bl_0_12
* pin bl_1_12
* pin br_1_12
* pin br_0_12
* pin bl_0_13
* pin bl_1_13
* pin br_1_13
* pin br_0_13
* pin bl_0_14
* pin bl_1_14
* pin br_1_14
* pin br_0_14
* pin bl_0_15
* pin bl_1_15
* pin br_1_15
* pin br_0_15
* pin bl_0_16
* pin bl_1_16
* pin br_1_16
* pin br_0_16
* pin bl_0_17
* pin bl_1_17
* pin br_1_17
* pin br_0_17
* pin bl_0_18
* pin bl_1_18
* pin br_1_18
* pin br_0_18
* pin bl_0_19
* pin bl_1_19
* pin br_1_19
* pin br_0_19
* pin bl_0_20
* pin bl_1_20
* pin br_1_20
* pin br_0_20
* pin bl_0_21
* pin bl_1_21
* pin br_1_21
* pin br_0_21
* pin bl_0_22
* pin bl_1_22
* pin br_1_22
* pin br_0_22
* pin bl_0_23
* pin bl_1_23
* pin br_1_23
* pin br_0_23
* pin bl_0_24
* pin bl_1_24
* pin br_1_24
* pin br_0_24
* pin bl_0_25
* pin bl_1_25
* pin br_1_25
* pin br_0_25
* pin bl_0_26
* pin bl_1_26
* pin br_1_26
* pin br_0_26
* pin bl_0_27
* pin bl_1_27
* pin br_1_27
* pin br_0_27
* pin bl_0_28
* pin bl_1_28
* pin br_1_28
* pin br_0_28
* pin bl_0_29
* pin bl_1_29
* pin br_1_29
* pin br_0_29
* pin bl_0_30
* pin bl_1_30
* pin br_1_30
* pin br_0_30
* pin bl_0_31
* pin bl_1_31
* pin br_1_31
* pin br_0_31
* pin rbl_bl_0_1
* pin rbl_bl_1_1
* pin rbl_br_1_1
* pin rbl_br_0_1
* pin wl_1_29
* pin wl_1_30
* pin wl_1_31
* pin wl_0_44
* pin wl_0_43
* pin wl_0_37
* pin wl_0_38
* pin wl_0_42
* pin wl_0_39
* pin wl_0_41
* pin wl_0_40
* pin wl_0_32
* pin wl_0_33
* pin wl_0_46
* pin wl_0_45
* pin wl_0_36
* pin wl_0_35
* pin wl_0_34
* pin wl_1_44
* pin wl_1_46
* pin wl_1_34
* pin wl_1_33
* pin wl_1_35
* pin wl_1_45
* pin wl_1_42
* pin wl_1_38
* pin wl_1_39
* pin wl_1_32
* pin wl_1_41
* pin wl_1_40
* pin wl_1_36
* pin wl_1_37
* pin wl_1_43
* pin wl_0_54
* pin wl_0_49
* pin wl_0_52
* pin wl_0_47
* pin wl_0_48
* pin wl_0_53
* pin wl_0_51
* pin wl_0_50
* pin wl_1_53
* pin wl_1_47
* pin wl_1_50
* pin wl_1_51
* pin wl_1_49
* pin wl_1_52
* pin wl_1_48
* pin wl_0_59
* pin wl_0_60
* pin wl_0_55
* pin wl_0_58
* pin wl_0_61
* pin wl_0_57
* pin wl_0_62
* pin wl_0_56
* pin wl_1_54
* pin wl_1_56
* pin wl_1_59
* pin wl_1_61
* pin wl_1_60
* pin wl_1_58
* pin wl_1_57
* pin wl_1_55
* pin wl_0_63
* pin rbl_wl_1_1
* pin wl_1_63
* pin wl_1_62
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_local_bitcell_array_1 1 2 3 4 5 6 7 8
+ 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 54 55 56 57 58 59 60 61 62 63 64
+ 65 66 67 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 114 115 116 117 118
+ 119 120 121 122 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139
+ 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158
+ 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177
+ 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196
+ 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215
+ 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234
+ 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250 251 252 253
+ 254 255 256 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275
+ 276 277 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322 323 324
+ 325 326 327 328 329 330 347 348 349 350 351 352 353 354 355 356 357 358 359
+ 360 361 377 378 379 380 381 382 383 384 385 390 391 392 393 394
* net 1 wl_0_3
* net 2 wl_0_4
* net 3 rbl_wl_0_0
* net 4 wl_0_1
* net 5 wl_0_0
* net 6 wl_0_6
* net 7 wl_0_2
* net 8 wl_0_5
* net 24 wl_1_1
* net 25 wl_1_0
* net 26 wl_1_6
* net 27 wl_1_2
* net 28 wl_1_4
* net 29 wl_1_3
* net 30 wl_1_5
* net 31 wl_0_9
* net 32 wl_0_10
* net 33 wl_0_8
* net 34 wl_0_11
* net 35 wl_0_12
* net 36 wl_0_7
* net 37 wl_0_13
* net 38 wl_0_14
* net 54 wl_1_7
* net 55 wl_1_13
* net 56 wl_1_8
* net 57 wl_1_9
* net 58 wl_1_10
* net 59 wl_1_11
* net 60 wl_1_12
* net 61 wl_0_20
* net 62 wl_0_17
* net 63 wl_0_16
* net 64 wl_0_18
* net 65 wl_0_19
* net 66 wl_0_15
* net 67 wl_0_21
* net 83 wl_1_15
* net 84 wl_1_14
* net 85 wl_1_21
* net 86 wl_1_18
* net 87 wl_1_19
* net 88 wl_1_17
* net 89 wl_1_16
* net 90 wl_1_20
* net 91 wl_0_27
* net 92 wl_0_24
* net 93 wl_0_28
* net 94 wl_0_23
* net 95 wl_0_29
* net 96 wl_0_22
* net 97 wl_0_26
* net 98 wl_0_25
* net 114 wl_1_24
* net 115 wl_1_22
* net 116 wl_1_27
* net 117 wl_1_28
* net 118 wl_1_25
* net 119 wl_1_26
* net 120 wl_1_23
* net 121 wl_0_30
* net 122 wl_0_31
* net 125 bl_0_0
* net 126 bl_1_0
* net 127 br_1_0
* net 128 br_0_0
* net 129 bl_0_1
* net 130 bl_1_1
* net 131 br_1_1
* net 132 br_0_1
* net 133 bl_0_2
* net 134 bl_1_2
* net 135 br_1_2
* net 136 br_0_2
* net 137 bl_0_3
* net 138 bl_1_3
* net 139 br_1_3
* net 140 br_0_3
* net 141 bl_0_4
* net 142 bl_1_4
* net 143 br_1_4
* net 144 br_0_4
* net 145 bl_0_5
* net 146 bl_1_5
* net 147 br_1_5
* net 148 br_0_5
* net 149 bl_0_6
* net 150 bl_1_6
* net 151 br_1_6
* net 152 br_0_6
* net 153 bl_0_7
* net 154 bl_1_7
* net 155 br_1_7
* net 156 br_0_7
* net 157 bl_0_8
* net 158 bl_1_8
* net 159 br_1_8
* net 160 br_0_8
* net 161 bl_0_9
* net 162 bl_1_9
* net 163 br_1_9
* net 164 br_0_9
* net 165 bl_0_10
* net 166 bl_1_10
* net 167 br_1_10
* net 168 br_0_10
* net 169 bl_0_11
* net 170 bl_1_11
* net 171 br_1_11
* net 172 br_0_11
* net 173 bl_0_12
* net 174 bl_1_12
* net 175 br_1_12
* net 176 br_0_12
* net 177 bl_0_13
* net 178 bl_1_13
* net 179 br_1_13
* net 180 br_0_13
* net 181 bl_0_14
* net 182 bl_1_14
* net 183 br_1_14
* net 184 br_0_14
* net 185 bl_0_15
* net 186 bl_1_15
* net 187 br_1_15
* net 188 br_0_15
* net 189 bl_0_16
* net 190 bl_1_16
* net 191 br_1_16
* net 192 br_0_16
* net 193 bl_0_17
* net 194 bl_1_17
* net 195 br_1_17
* net 196 br_0_17
* net 197 bl_0_18
* net 198 bl_1_18
* net 199 br_1_18
* net 200 br_0_18
* net 201 bl_0_19
* net 202 bl_1_19
* net 203 br_1_19
* net 204 br_0_19
* net 205 bl_0_20
* net 206 bl_1_20
* net 207 br_1_20
* net 208 br_0_20
* net 209 bl_0_21
* net 210 bl_1_21
* net 211 br_1_21
* net 212 br_0_21
* net 213 bl_0_22
* net 214 bl_1_22
* net 215 br_1_22
* net 216 br_0_22
* net 217 bl_0_23
* net 218 bl_1_23
* net 219 br_1_23
* net 220 br_0_23
* net 221 bl_0_24
* net 222 bl_1_24
* net 223 br_1_24
* net 224 br_0_24
* net 225 bl_0_25
* net 226 bl_1_25
* net 227 br_1_25
* net 228 br_0_25
* net 229 bl_0_26
* net 230 bl_1_26
* net 231 br_1_26
* net 232 br_0_26
* net 233 bl_0_27
* net 234 bl_1_27
* net 235 br_1_27
* net 236 br_0_27
* net 237 bl_0_28
* net 238 bl_1_28
* net 239 br_1_28
* net 240 br_0_28
* net 241 bl_0_29
* net 242 bl_1_29
* net 243 br_1_29
* net 244 br_0_29
* net 245 bl_0_30
* net 246 bl_1_30
* net 247 br_1_30
* net 248 br_0_30
* net 249 bl_0_31
* net 250 bl_1_31
* net 251 br_1_31
* net 252 br_0_31
* net 253 rbl_bl_0_1
* net 254 rbl_bl_1_1
* net 255 rbl_br_1_1
* net 256 rbl_br_0_1
* net 260 wl_1_29
* net 261 wl_1_30
* net 262 wl_1_31
* net 263 wl_0_44
* net 264 wl_0_43
* net 265 wl_0_37
* net 266 wl_0_38
* net 267 wl_0_42
* net 268 wl_0_39
* net 269 wl_0_41
* net 270 wl_0_40
* net 271 wl_0_32
* net 272 wl_0_33
* net 273 wl_0_46
* net 274 wl_0_45
* net 275 wl_0_36
* net 276 wl_0_35
* net 277 wl_0_34
* net 308 wl_1_44
* net 309 wl_1_46
* net 310 wl_1_34
* net 311 wl_1_33
* net 312 wl_1_35
* net 313 wl_1_45
* net 314 wl_1_42
* net 315 wl_1_38
* net 316 wl_1_39
* net 317 wl_1_32
* net 318 wl_1_41
* net 319 wl_1_40
* net 320 wl_1_36
* net 321 wl_1_37
* net 322 wl_1_43
* net 323 wl_0_54
* net 324 wl_0_49
* net 325 wl_0_52
* net 326 wl_0_47
* net 327 wl_0_48
* net 328 wl_0_53
* net 329 wl_0_51
* net 330 wl_0_50
* net 347 wl_1_53
* net 348 wl_1_47
* net 349 wl_1_50
* net 350 wl_1_51
* net 351 wl_1_49
* net 352 wl_1_52
* net 353 wl_1_48
* net 354 wl_0_59
* net 355 wl_0_60
* net 356 wl_0_55
* net 357 wl_0_58
* net 358 wl_0_61
* net 359 wl_0_57
* net 360 wl_0_62
* net 361 wl_0_56
* net 377 wl_1_54
* net 378 wl_1_56
* net 379 wl_1_59
* net 380 wl_1_61
* net 381 wl_1_60
* net 382 wl_1_58
* net 383 wl_1_57
* net 384 wl_1_55
* net 385 wl_0_63
* net 390 rbl_wl_1_1
* net 391 wl_1_63
* net 392 wl_1_62
* net 393 vdd
* net 394 gnd
* cell instance $3 r0 *1 0,1.745
X$3 3 11 5 10 4 9 7 12 1 16 2 15 8 14 6 13 36 41 33 39 31 45 32 40 34 42 35 44
+ 37 43 38 71 66 68 63 75 62 74 64 69 65 70 61 73 67 72 96 101 94 102 92 103 98
+ 105 97 99 91 104 93 106 95 100 121 124 122 123 271 278 272 282 277 281 276
+ 280 275 285 265 291 266 290 268 288 270 286 269 287 267 289 264 292 263 279
+ 274 283 273 284 326 331 327 338 324 334 330 335 329 336 325 332 328 333 323
+ 337 356 362 361 363 359 368 357 367 354 366 355 365 358 364 360 387 385 386
+ 393 394 custom_sram_1r1w_32_256_freepdk45_wordline_buffer_array
* cell instance $18 r0 *1 6.3325,0
X$18 52 102 11 75 74 76 107 45 69 108 81 103 70 73 46 49 71 50 43 44 48 82 68
+ 79 101 42 40 72 53 78 77 80 112 39 19 10 9 21 22 12 16 23 20 15 14 51 47 41
+ 13 17 18 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179
+ 180 181 182 183 184 185 186 187 188 189 190 258 257 124 123 100 106 110 109
+ 104 105 99 259 111 113 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 331 340 388 345
+ 376 343 284 363 297 332 283 334 333 282 339 335 346 342 336 341 344 337 365
+ 305 338 362 372 281 370 374 369 298 366 306 387 285 295 296 287 278 371 286
+ 307 367 304 288 291 300 290 301 302 364 375 289 279 294 280 293 389 292 299
+ 373 368 386 303 393 394
+ custom_sram_1r1w_32_256_freepdk45_capped_replica_bitcell_array_1
* cell instance $19 r180 *1 55.66,100.415
X$19 390 388 391 389 392 371 380 373 381 370 379 369 382 375 383 374 378 376
+ 384 372 377 342 347 339 352 340 350 345 349 346 351 341 353 343 348 344 309
+ 297 313 296 308 294 322 293 314 298 318 295 319 307 316 304 315 301 321 300
+ 320 306 312 303 310 305 311 299 317 302 262 258 261 257 260 259 117 110 116
+ 109 119 111 118 113 114 108 120 107 115 112 85 78 90 77 87 76 86 82 88 81 89
+ 80 83 79 84 49 55 50 60 48 59 46 58 53 57 52 56 51 54 47 26 17 30 18 28 20 29
+ 23 27 22 24 21 25 19 393 394
+ custom_sram_1r1w_32_256_freepdk45_wordline_buffer_array
.ENDS custom_sram_1r1w_32_256_freepdk45_local_bitcell_array_1

* cell custom_sram_1r1w_32_256_freepdk45_local_bitcell_array_0
* pin wl_0_1
* pin wl_0_2
* pin wl_0_3
* pin wl_0_4
* pin wl_0_0
* pin rbl_wl_0_0
* pin wl_0_6
* pin wl_0_5
* pin wl_1_5
* pin wl_1_1
* pin wl_1_3
* pin wl_1_0
* pin wl_1_2
* pin wl_1_4
* pin wl_0_13
* pin wl_0_9
* pin wl_0_12
* pin wl_0_10
* pin wl_0_8
* pin wl_0_7
* pin wl_0_11
* pin wl_1_6
* pin wl_1_7
* pin wl_1_13
* pin wl_1_10
* pin wl_1_11
* pin wl_1_9
* pin wl_1_8
* pin wl_1_12
* pin wl_0_17
* pin wl_0_18
* pin wl_0_16
* pin wl_0_15
* pin wl_0_19
* pin wl_0_21
* pin wl_0_14
* pin wl_0_20
* pin wl_1_15
* pin wl_1_20
* pin wl_1_14
* pin wl_1_19
* pin wl_1_16
* pin wl_1_17
* pin wl_1_18
* pin wl_0_24
* pin wl_0_23
* pin wl_0_25
* pin wl_0_26
* pin wl_0_22
* pin wl_0_27
* pin wl_0_28
* pin wl_1_28
* pin wl_1_27
* pin wl_1_21
* pin wl_1_24
* pin wl_1_25
* pin wl_1_23
* pin wl_1_26
* pin wl_1_22
* pin wl_0_30
* pin wl_0_29
* pin wl_0_31
* pin bl_0_0
* pin bl_1_0
* pin br_1_0
* pin br_0_0
* pin bl_0_1
* pin bl_1_1
* pin br_1_1
* pin br_0_1
* pin bl_0_2
* pin bl_1_2
* pin br_1_2
* pin br_0_2
* pin bl_0_3
* pin bl_1_3
* pin br_1_3
* pin br_0_3
* pin bl_0_4
* pin bl_1_4
* pin br_1_4
* pin br_0_4
* pin bl_0_5
* pin bl_1_5
* pin br_1_5
* pin br_0_5
* pin bl_0_6
* pin bl_1_6
* pin br_1_6
* pin br_0_6
* pin bl_0_7
* pin bl_1_7
* pin br_1_7
* pin br_0_7
* pin bl_0_8
* pin bl_1_8
* pin br_1_8
* pin br_0_8
* pin bl_0_9
* pin bl_1_9
* pin br_1_9
* pin br_0_9
* pin bl_0_10
* pin bl_1_10
* pin br_1_10
* pin br_0_10
* pin bl_0_11
* pin bl_1_11
* pin br_1_11
* pin br_0_11
* pin bl_0_12
* pin bl_1_12
* pin br_1_12
* pin br_0_12
* pin bl_0_13
* pin bl_1_13
* pin br_1_13
* pin br_0_13
* pin bl_0_14
* pin bl_1_14
* pin br_1_14
* pin br_0_14
* pin bl_0_15
* pin bl_1_15
* pin br_1_15
* pin br_0_15
* pin bl_0_16
* pin bl_1_16
* pin br_1_16
* pin br_0_16
* pin bl_0_17
* pin bl_1_17
* pin br_1_17
* pin br_0_17
* pin bl_0_18
* pin bl_1_18
* pin br_1_18
* pin br_0_18
* pin bl_0_19
* pin bl_1_19
* pin br_1_19
* pin br_0_19
* pin bl_0_20
* pin bl_1_20
* pin br_1_20
* pin br_0_20
* pin bl_0_21
* pin bl_1_21
* pin br_1_21
* pin br_0_21
* pin bl_0_22
* pin bl_1_22
* pin br_1_22
* pin br_0_22
* pin bl_0_23
* pin bl_1_23
* pin br_1_23
* pin br_0_23
* pin bl_0_24
* pin bl_1_24
* pin br_1_24
* pin br_0_24
* pin bl_0_25
* pin bl_1_25
* pin br_1_25
* pin br_0_25
* pin bl_0_26
* pin bl_1_26
* pin br_1_26
* pin br_0_26
* pin bl_0_27
* pin bl_1_27
* pin br_1_27
* pin br_0_27
* pin bl_0_28
* pin bl_1_28
* pin br_1_28
* pin br_0_28
* pin bl_0_29
* pin bl_1_29
* pin br_1_29
* pin br_0_29
* pin bl_0_30
* pin bl_1_30
* pin br_1_30
* pin br_0_30
* pin bl_0_31
* pin bl_1_31
* pin br_1_31
* pin br_0_31
* pin wl_1_31
* pin wl_1_29
* pin wl_1_30
* pin wl_0_37
* pin wl_0_34
* pin wl_0_38
* pin wl_0_39
* pin wl_0_35
* pin wl_0_40
* pin wl_0_42
* pin wl_0_41
* pin wl_0_32
* pin wl_0_33
* pin wl_0_36
* pin wl_0_46
* pin wl_0_45
* pin wl_0_43
* pin wl_0_44
* pin wl_1_34
* pin wl_1_40
* pin wl_1_45
* pin wl_1_39
* pin wl_1_38
* pin wl_1_35
* pin wl_1_32
* pin wl_1_33
* pin wl_1_43
* pin wl_1_42
* pin wl_1_37
* pin wl_1_44
* pin wl_1_36
* pin wl_1_41
* pin wl_0_53
* pin wl_0_47
* pin wl_0_52
* pin wl_0_48
* pin wl_0_51
* pin wl_0_50
* pin wl_0_49
* pin wl_1_48
* pin wl_1_53
* pin wl_1_51
* pin wl_1_46
* pin wl_1_50
* pin wl_1_52
* pin wl_1_47
* pin wl_1_49
* pin wl_0_57
* pin wl_0_58
* pin wl_0_55
* pin wl_0_56
* pin wl_0_59
* pin wl_0_60
* pin wl_0_61
* pin wl_0_54
* pin wl_1_55
* pin wl_1_60
* pin wl_1_54
* pin wl_1_59
* pin wl_1_56
* pin wl_1_57
* pin wl_1_58
* pin wl_0_62
* pin wl_0_63
* pin rbl_wl_1_1
* pin wl_1_61
* pin wl_1_63
* pin wl_1_62
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_local_bitcell_array_0 1 2 3 4 5 6 7 8
+ 24 25 26 27 28 29 30 31 32 33 34 35 36 52 53 54 55 56 57 58 59 60 61 62 63 64
+ 65 66 67 82 83 84 85 86 87 88 89 90 91 92 93 94 95 111 112 113 114 115 116
+ 117 118 119 120 121 125 126 127 128 129 130 131 132 133 134 135 136 137 138
+ 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157
+ 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176
+ 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195
+ 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214
+ 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233
+ 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250 251 252
+ 256 257 258 259 260 261 262 263 264 265 266 267 268 269 270 271 272 273 304
+ 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322 323
+ 324 340 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 370 371
+ 372 373 374 375 376 377 378 385 386 387 388 389 390
* net 1 wl_0_1
* net 2 wl_0_2
* net 3 wl_0_3
* net 4 wl_0_4
* net 5 wl_0_0
* net 6 rbl_wl_0_0
* net 7 wl_0_6
* net 8 wl_0_5
* net 24 wl_1_5
* net 25 wl_1_1
* net 26 wl_1_3
* net 27 wl_1_0
* net 28 wl_1_2
* net 29 wl_1_4
* net 30 wl_0_13
* net 31 wl_0_9
* net 32 wl_0_12
* net 33 wl_0_10
* net 34 wl_0_8
* net 35 wl_0_7
* net 36 wl_0_11
* net 52 wl_1_6
* net 53 wl_1_7
* net 54 wl_1_13
* net 55 wl_1_10
* net 56 wl_1_11
* net 57 wl_1_9
* net 58 wl_1_8
* net 59 wl_1_12
* net 60 wl_0_17
* net 61 wl_0_18
* net 62 wl_0_16
* net 63 wl_0_15
* net 64 wl_0_19
* net 65 wl_0_21
* net 66 wl_0_14
* net 67 wl_0_20
* net 82 wl_1_15
* net 83 wl_1_20
* net 84 wl_1_14
* net 85 wl_1_19
* net 86 wl_1_16
* net 87 wl_1_17
* net 88 wl_1_18
* net 89 wl_0_24
* net 90 wl_0_23
* net 91 wl_0_25
* net 92 wl_0_26
* net 93 wl_0_22
* net 94 wl_0_27
* net 95 wl_0_28
* net 111 wl_1_28
* net 112 wl_1_27
* net 113 wl_1_21
* net 114 wl_1_24
* net 115 wl_1_25
* net 116 wl_1_23
* net 117 wl_1_26
* net 118 wl_1_22
* net 119 wl_0_30
* net 120 wl_0_29
* net 121 wl_0_31
* net 125 bl_0_0
* net 126 bl_1_0
* net 127 br_1_0
* net 128 br_0_0
* net 129 bl_0_1
* net 130 bl_1_1
* net 131 br_1_1
* net 132 br_0_1
* net 133 bl_0_2
* net 134 bl_1_2
* net 135 br_1_2
* net 136 br_0_2
* net 137 bl_0_3
* net 138 bl_1_3
* net 139 br_1_3
* net 140 br_0_3
* net 141 bl_0_4
* net 142 bl_1_4
* net 143 br_1_4
* net 144 br_0_4
* net 145 bl_0_5
* net 146 bl_1_5
* net 147 br_1_5
* net 148 br_0_5
* net 149 bl_0_6
* net 150 bl_1_6
* net 151 br_1_6
* net 152 br_0_6
* net 153 bl_0_7
* net 154 bl_1_7
* net 155 br_1_7
* net 156 br_0_7
* net 157 bl_0_8
* net 158 bl_1_8
* net 159 br_1_8
* net 160 br_0_8
* net 161 bl_0_9
* net 162 bl_1_9
* net 163 br_1_9
* net 164 br_0_9
* net 165 bl_0_10
* net 166 bl_1_10
* net 167 br_1_10
* net 168 br_0_10
* net 169 bl_0_11
* net 170 bl_1_11
* net 171 br_1_11
* net 172 br_0_11
* net 173 bl_0_12
* net 174 bl_1_12
* net 175 br_1_12
* net 176 br_0_12
* net 177 bl_0_13
* net 178 bl_1_13
* net 179 br_1_13
* net 180 br_0_13
* net 181 bl_0_14
* net 182 bl_1_14
* net 183 br_1_14
* net 184 br_0_14
* net 185 bl_0_15
* net 186 bl_1_15
* net 187 br_1_15
* net 188 br_0_15
* net 189 bl_0_16
* net 190 bl_1_16
* net 191 br_1_16
* net 192 br_0_16
* net 193 bl_0_17
* net 194 bl_1_17
* net 195 br_1_17
* net 196 br_0_17
* net 197 bl_0_18
* net 198 bl_1_18
* net 199 br_1_18
* net 200 br_0_18
* net 201 bl_0_19
* net 202 bl_1_19
* net 203 br_1_19
* net 204 br_0_19
* net 205 bl_0_20
* net 206 bl_1_20
* net 207 br_1_20
* net 208 br_0_20
* net 209 bl_0_21
* net 210 bl_1_21
* net 211 br_1_21
* net 212 br_0_21
* net 213 bl_0_22
* net 214 bl_1_22
* net 215 br_1_22
* net 216 br_0_22
* net 217 bl_0_23
* net 218 bl_1_23
* net 219 br_1_23
* net 220 br_0_23
* net 221 bl_0_24
* net 222 bl_1_24
* net 223 br_1_24
* net 224 br_0_24
* net 225 bl_0_25
* net 226 bl_1_25
* net 227 br_1_25
* net 228 br_0_25
* net 229 bl_0_26
* net 230 bl_1_26
* net 231 br_1_26
* net 232 br_0_26
* net 233 bl_0_27
* net 234 bl_1_27
* net 235 br_1_27
* net 236 br_0_27
* net 237 bl_0_28
* net 238 bl_1_28
* net 239 br_1_28
* net 240 br_0_28
* net 241 bl_0_29
* net 242 bl_1_29
* net 243 br_1_29
* net 244 br_0_29
* net 245 bl_0_30
* net 246 bl_1_30
* net 247 br_1_30
* net 248 br_0_30
* net 249 bl_0_31
* net 250 bl_1_31
* net 251 br_1_31
* net 252 br_0_31
* net 256 wl_1_31
* net 257 wl_1_29
* net 258 wl_1_30
* net 259 wl_0_37
* net 260 wl_0_34
* net 261 wl_0_38
* net 262 wl_0_39
* net 263 wl_0_35
* net 264 wl_0_40
* net 265 wl_0_42
* net 266 wl_0_41
* net 267 wl_0_32
* net 268 wl_0_33
* net 269 wl_0_36
* net 270 wl_0_46
* net 271 wl_0_45
* net 272 wl_0_43
* net 273 wl_0_44
* net 304 wl_1_34
* net 305 wl_1_40
* net 306 wl_1_45
* net 307 wl_1_39
* net 308 wl_1_38
* net 309 wl_1_35
* net 310 wl_1_32
* net 311 wl_1_33
* net 312 wl_1_43
* net 313 wl_1_42
* net 314 wl_1_37
* net 315 wl_1_44
* net 316 wl_1_36
* net 317 wl_1_41
* net 318 wl_0_53
* net 319 wl_0_47
* net 320 wl_0_52
* net 321 wl_0_48
* net 322 wl_0_51
* net 323 wl_0_50
* net 324 wl_0_49
* net 340 wl_1_48
* net 341 wl_1_53
* net 342 wl_1_51
* net 343 wl_1_46
* net 344 wl_1_50
* net 345 wl_1_52
* net 346 wl_1_47
* net 347 wl_1_49
* net 348 wl_0_57
* net 349 wl_0_58
* net 350 wl_0_55
* net 351 wl_0_56
* net 352 wl_0_59
* net 353 wl_0_60
* net 354 wl_0_61
* net 355 wl_0_54
* net 370 wl_1_55
* net 371 wl_1_60
* net 372 wl_1_54
* net 373 wl_1_59
* net 374 wl_1_56
* net 375 wl_1_57
* net 376 wl_1_58
* net 377 wl_0_62
* net 378 wl_0_63
* net 385 rbl_wl_1_1
* net 386 wl_1_61
* net 387 wl_1_63
* net 388 wl_1_62
* net 389 vdd
* net 390 gnd
* cell instance $3 r0 *1 0,1.745
X$3 6 11 5 10 1 9 2 12 3 16 4 15 8 14 7 13 35 37 34 43 31 41 33 40 36 39 32 42
+ 30 38 66 70 63 69 62 68 60 75 61 74 64 72 67 71 65 73 93 96 90 97 89 102 91
+ 101 92 98 94 100 95 99 120 124 119 122 121 123 267 284 268 280 260 278 263
+ 275 269 287 259 286 261 279 262 285 264 282 266 277 265 283 272 276 273 281
+ 271 274 270 288 319 327 321 331 324 325 323 328 322 329 320 330 318 326 355
+ 357 350 358 351 356 348 363 349 362 352 361 353 360 354 359 377 380 378 379
+ 389 390 custom_sram_1r1w_32_256_freepdk45_wordline_buffer_array
* cell instance $18 r0 *1 6.3325,0
X$18 48 79 76 41 107 72 43 74 49 80 47 42 97 22 51 71 40 73 77 96 39 105 46 108
+ 17 78 18 19 14 10 9 20 70 69 15 12 21 44 16 38 68 50 45 37 23 11 13 75 81 125
+ 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144
+ 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 100 122 253 109 254 102 124 101 123 110 255 104 99 98
+ 106 103 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205
+ 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224
+ 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243
+ 244 245 246 247 248 249 250 251 252 384 380 382 339 325 331 335 379 338 381
+ 336 328 327 361 366 362 365 368 284 369 363 364 356 367 360 329 358 359 357
+ 332 337 326 330 334 333 383 285 281 275 297 303 294 287 286 292 290 279 288
+ 300 293 302 282 276 277 295 296 283 274 278 289 291 301 280 299 298 389 390
+ custom_sram_1r1w_32_256_freepdk45_capped_replica_bitcell_array_0
* cell instance $19 r180 *1 54.485,100.415
X$19 385 382 387 381 388 384 386 383 371 364 373 368 376 365 375 369 374 367
+ 370 366 372 332 341 337 345 334 342 333 344 338 347 339 340 335 346 336 343
+ 298 306 301 315 294 312 293 313 296 317 295 305 302 307 300 308 290 314 292
+ 316 303 309 297 304 289 311 291 310 299 256 255 258 253 257 254 111 106 112
+ 103 117 104 115 110 114 109 116 107 118 108 113 105 83 79 85 76 88 80 87 81
+ 86 78 82 77 84 45 54 44 59 47 56 46 55 51 57 48 58 49 53 50 52 23 24 18 29 21
+ 26 22 28 17 25 20 27 19 389 390
+ custom_sram_1r1w_32_256_freepdk45_wordline_buffer_array
.ENDS custom_sram_1r1w_32_256_freepdk45_local_bitcell_array_0

* cell custom_sram_1r1w_32_256_freepdk45_local_bitcell_array
* pin wl_0_3
* pin wl_0_4
* pin rbl_wl_0_0
* pin wl_0_1
* pin wl_0_0
* pin wl_0_6
* pin wl_0_2
* pin wl_0_5
* pin wl_1_1
* pin wl_1_0
* pin wl_1_6
* pin wl_1_2
* pin wl_1_4
* pin wl_1_3
* pin wl_1_5
* pin wl_0_9
* pin wl_0_10
* pin wl_0_8
* pin wl_0_11
* pin wl_0_12
* pin wl_0_7
* pin wl_0_13
* pin wl_0_14
* pin wl_1_7
* pin wl_1_13
* pin wl_1_8
* pin wl_1_9
* pin wl_1_10
* pin wl_1_11
* pin wl_1_12
* pin wl_0_20
* pin wl_0_17
* pin wl_0_16
* pin wl_0_18
* pin wl_0_19
* pin wl_0_15
* pin wl_0_21
* pin wl_1_15
* pin wl_1_14
* pin wl_1_21
* pin wl_1_18
* pin wl_1_19
* pin wl_1_17
* pin wl_1_16
* pin wl_1_20
* pin wl_0_27
* pin wl_0_24
* pin wl_0_28
* pin wl_0_23
* pin wl_0_29
* pin wl_0_22
* pin wl_0_26
* pin wl_0_25
* pin wl_1_24
* pin wl_1_22
* pin wl_1_27
* pin wl_1_28
* pin wl_1_25
* pin wl_1_26
* pin wl_1_23
* pin wl_0_30
* pin wl_0_31
* pin rbl_bl_0_0
* pin rbl_bl_1_0
* pin rbl_br_1_0
* pin rbl_br_0_0
* pin bl_0_0
* pin bl_1_0
* pin br_1_0
* pin br_0_0
* pin bl_0_1
* pin bl_1_1
* pin br_1_1
* pin br_0_1
* pin bl_0_2
* pin bl_1_2
* pin br_1_2
* pin br_0_2
* pin bl_0_3
* pin bl_1_3
* pin br_1_3
* pin br_0_3
* pin bl_0_4
* pin bl_1_4
* pin br_1_4
* pin br_0_4
* pin bl_0_5
* pin bl_1_5
* pin br_1_5
* pin br_0_5
* pin bl_0_6
* pin bl_1_6
* pin br_1_6
* pin br_0_6
* pin bl_0_7
* pin bl_1_7
* pin br_1_7
* pin br_0_7
* pin bl_0_8
* pin bl_1_8
* pin br_1_8
* pin br_0_8
* pin bl_0_9
* pin bl_1_9
* pin br_1_9
* pin br_0_9
* pin bl_0_10
* pin bl_1_10
* pin br_1_10
* pin br_0_10
* pin bl_0_11
* pin bl_1_11
* pin br_1_11
* pin br_0_11
* pin bl_0_12
* pin bl_1_12
* pin br_1_12
* pin br_0_12
* pin bl_0_13
* pin bl_1_13
* pin br_1_13
* pin br_0_13
* pin bl_0_14
* pin bl_1_14
* pin br_1_14
* pin br_0_14
* pin bl_0_15
* pin bl_1_15
* pin br_1_15
* pin br_0_15
* pin bl_0_16
* pin bl_1_16
* pin br_1_16
* pin br_0_16
* pin bl_0_17
* pin bl_1_17
* pin br_1_17
* pin br_0_17
* pin bl_0_18
* pin bl_1_18
* pin br_1_18
* pin br_0_18
* pin bl_0_19
* pin bl_1_19
* pin br_1_19
* pin br_0_19
* pin bl_0_20
* pin bl_1_20
* pin br_1_20
* pin br_0_20
* pin bl_0_21
* pin bl_1_21
* pin br_1_21
* pin br_0_21
* pin bl_0_22
* pin bl_1_22
* pin br_1_22
* pin br_0_22
* pin bl_0_23
* pin bl_1_23
* pin br_1_23
* pin br_0_23
* pin bl_0_24
* pin bl_1_24
* pin br_1_24
* pin br_0_24
* pin bl_0_25
* pin bl_1_25
* pin br_1_25
* pin br_0_25
* pin bl_0_26
* pin bl_1_26
* pin br_1_26
* pin br_0_26
* pin bl_0_27
* pin bl_1_27
* pin br_1_27
* pin br_0_27
* pin bl_0_28
* pin bl_1_28
* pin br_1_28
* pin br_0_28
* pin bl_0_29
* pin bl_1_29
* pin br_1_29
* pin br_0_29
* pin bl_0_30
* pin bl_1_30
* pin br_1_30
* pin br_0_30
* pin bl_0_31
* pin bl_1_31
* pin br_1_31
* pin br_0_31
* pin wl_1_29
* pin wl_1_30
* pin wl_1_31
* pin wl_0_44
* pin wl_0_43
* pin wl_0_37
* pin wl_0_38
* pin wl_0_42
* pin wl_0_39
* pin wl_0_41
* pin wl_0_40
* pin wl_0_32
* pin wl_0_33
* pin wl_0_46
* pin wl_0_45
* pin wl_0_36
* pin wl_0_35
* pin wl_0_34
* pin wl_1_44
* pin wl_1_46
* pin wl_1_34
* pin wl_1_33
* pin wl_1_35
* pin wl_1_45
* pin wl_1_42
* pin wl_1_38
* pin wl_1_39
* pin wl_1_32
* pin wl_1_41
* pin wl_1_40
* pin wl_1_36
* pin wl_1_37
* pin wl_1_43
* pin wl_0_54
* pin wl_0_49
* pin wl_0_52
* pin wl_0_47
* pin wl_0_48
* pin wl_0_53
* pin wl_0_51
* pin wl_0_50
* pin wl_1_53
* pin wl_1_47
* pin wl_1_50
* pin wl_1_51
* pin wl_1_49
* pin wl_1_52
* pin wl_1_48
* pin wl_0_59
* pin wl_0_60
* pin wl_0_55
* pin wl_0_58
* pin wl_0_61
* pin wl_0_57
* pin wl_0_62
* pin wl_0_56
* pin wl_1_54
* pin wl_1_56
* pin wl_1_59
* pin wl_1_61
* pin wl_1_60
* pin wl_1_58
* pin wl_1_57
* pin wl_1_55
* pin wl_0_63
* pin rbl_wl_1_1
* pin wl_1_63
* pin wl_1_62
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_local_bitcell_array 1 2 3 4 5 6 7 8
+ 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 54 55 56 57 58 59 60 61 62 63 64
+ 65 66 67 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 114 115 116 117 118
+ 119 120 121 122 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139
+ 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158
+ 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177
+ 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196
+ 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215
+ 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234
+ 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250 251 252 253
+ 254 255 256 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275
+ 276 277 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322 323 324
+ 325 326 327 328 329 330 347 348 349 350 351 352 353 354 355 356 357 358 359
+ 360 361 377 378 379 380 381 382 383 384 385 390 391 392 393 394
* net 1 wl_0_3
* net 2 wl_0_4
* net 3 rbl_wl_0_0
* net 4 wl_0_1
* net 5 wl_0_0
* net 6 wl_0_6
* net 7 wl_0_2
* net 8 wl_0_5
* net 24 wl_1_1
* net 25 wl_1_0
* net 26 wl_1_6
* net 27 wl_1_2
* net 28 wl_1_4
* net 29 wl_1_3
* net 30 wl_1_5
* net 31 wl_0_9
* net 32 wl_0_10
* net 33 wl_0_8
* net 34 wl_0_11
* net 35 wl_0_12
* net 36 wl_0_7
* net 37 wl_0_13
* net 38 wl_0_14
* net 54 wl_1_7
* net 55 wl_1_13
* net 56 wl_1_8
* net 57 wl_1_9
* net 58 wl_1_10
* net 59 wl_1_11
* net 60 wl_1_12
* net 61 wl_0_20
* net 62 wl_0_17
* net 63 wl_0_16
* net 64 wl_0_18
* net 65 wl_0_19
* net 66 wl_0_15
* net 67 wl_0_21
* net 83 wl_1_15
* net 84 wl_1_14
* net 85 wl_1_21
* net 86 wl_1_18
* net 87 wl_1_19
* net 88 wl_1_17
* net 89 wl_1_16
* net 90 wl_1_20
* net 91 wl_0_27
* net 92 wl_0_24
* net 93 wl_0_28
* net 94 wl_0_23
* net 95 wl_0_29
* net 96 wl_0_22
* net 97 wl_0_26
* net 98 wl_0_25
* net 114 wl_1_24
* net 115 wl_1_22
* net 116 wl_1_27
* net 117 wl_1_28
* net 118 wl_1_25
* net 119 wl_1_26
* net 120 wl_1_23
* net 121 wl_0_30
* net 122 wl_0_31
* net 125 rbl_bl_0_0
* net 126 rbl_bl_1_0
* net 127 rbl_br_1_0
* net 128 rbl_br_0_0
* net 129 bl_0_0
* net 130 bl_1_0
* net 131 br_1_0
* net 132 br_0_0
* net 133 bl_0_1
* net 134 bl_1_1
* net 135 br_1_1
* net 136 br_0_1
* net 137 bl_0_2
* net 138 bl_1_2
* net 139 br_1_2
* net 140 br_0_2
* net 141 bl_0_3
* net 142 bl_1_3
* net 143 br_1_3
* net 144 br_0_3
* net 145 bl_0_4
* net 146 bl_1_4
* net 147 br_1_4
* net 148 br_0_4
* net 149 bl_0_5
* net 150 bl_1_5
* net 151 br_1_5
* net 152 br_0_5
* net 153 bl_0_6
* net 154 bl_1_6
* net 155 br_1_6
* net 156 br_0_6
* net 157 bl_0_7
* net 158 bl_1_7
* net 159 br_1_7
* net 160 br_0_7
* net 161 bl_0_8
* net 162 bl_1_8
* net 163 br_1_8
* net 164 br_0_8
* net 165 bl_0_9
* net 166 bl_1_9
* net 167 br_1_9
* net 168 br_0_9
* net 169 bl_0_10
* net 170 bl_1_10
* net 171 br_1_10
* net 172 br_0_10
* net 173 bl_0_11
* net 174 bl_1_11
* net 175 br_1_11
* net 176 br_0_11
* net 177 bl_0_12
* net 178 bl_1_12
* net 179 br_1_12
* net 180 br_0_12
* net 181 bl_0_13
* net 182 bl_1_13
* net 183 br_1_13
* net 184 br_0_13
* net 185 bl_0_14
* net 186 bl_1_14
* net 187 br_1_14
* net 188 br_0_14
* net 189 bl_0_15
* net 190 bl_1_15
* net 191 br_1_15
* net 192 br_0_15
* net 193 bl_0_16
* net 194 bl_1_16
* net 195 br_1_16
* net 196 br_0_16
* net 197 bl_0_17
* net 198 bl_1_17
* net 199 br_1_17
* net 200 br_0_17
* net 201 bl_0_18
* net 202 bl_1_18
* net 203 br_1_18
* net 204 br_0_18
* net 205 bl_0_19
* net 206 bl_1_19
* net 207 br_1_19
* net 208 br_0_19
* net 209 bl_0_20
* net 210 bl_1_20
* net 211 br_1_20
* net 212 br_0_20
* net 213 bl_0_21
* net 214 bl_1_21
* net 215 br_1_21
* net 216 br_0_21
* net 217 bl_0_22
* net 218 bl_1_22
* net 219 br_1_22
* net 220 br_0_22
* net 221 bl_0_23
* net 222 bl_1_23
* net 223 br_1_23
* net 224 br_0_23
* net 225 bl_0_24
* net 226 bl_1_24
* net 227 br_1_24
* net 228 br_0_24
* net 229 bl_0_25
* net 230 bl_1_25
* net 231 br_1_25
* net 232 br_0_25
* net 233 bl_0_26
* net 234 bl_1_26
* net 235 br_1_26
* net 236 br_0_26
* net 237 bl_0_27
* net 238 bl_1_27
* net 239 br_1_27
* net 240 br_0_27
* net 241 bl_0_28
* net 242 bl_1_28
* net 243 br_1_28
* net 244 br_0_28
* net 245 bl_0_29
* net 246 bl_1_29
* net 247 br_1_29
* net 248 br_0_29
* net 249 bl_0_30
* net 250 bl_1_30
* net 251 br_1_30
* net 252 br_0_30
* net 253 bl_0_31
* net 254 bl_1_31
* net 255 br_1_31
* net 256 br_0_31
* net 260 wl_1_29
* net 261 wl_1_30
* net 262 wl_1_31
* net 263 wl_0_44
* net 264 wl_0_43
* net 265 wl_0_37
* net 266 wl_0_38
* net 267 wl_0_42
* net 268 wl_0_39
* net 269 wl_0_41
* net 270 wl_0_40
* net 271 wl_0_32
* net 272 wl_0_33
* net 273 wl_0_46
* net 274 wl_0_45
* net 275 wl_0_36
* net 276 wl_0_35
* net 277 wl_0_34
* net 308 wl_1_44
* net 309 wl_1_46
* net 310 wl_1_34
* net 311 wl_1_33
* net 312 wl_1_35
* net 313 wl_1_45
* net 314 wl_1_42
* net 315 wl_1_38
* net 316 wl_1_39
* net 317 wl_1_32
* net 318 wl_1_41
* net 319 wl_1_40
* net 320 wl_1_36
* net 321 wl_1_37
* net 322 wl_1_43
* net 323 wl_0_54
* net 324 wl_0_49
* net 325 wl_0_52
* net 326 wl_0_47
* net 327 wl_0_48
* net 328 wl_0_53
* net 329 wl_0_51
* net 330 wl_0_50
* net 347 wl_1_53
* net 348 wl_1_47
* net 349 wl_1_50
* net 350 wl_1_51
* net 351 wl_1_49
* net 352 wl_1_52
* net 353 wl_1_48
* net 354 wl_0_59
* net 355 wl_0_60
* net 356 wl_0_55
* net 357 wl_0_58
* net 358 wl_0_61
* net 359 wl_0_57
* net 360 wl_0_62
* net 361 wl_0_56
* net 377 wl_1_54
* net 378 wl_1_56
* net 379 wl_1_59
* net 380 wl_1_61
* net 381 wl_1_60
* net 382 wl_1_58
* net 383 wl_1_57
* net 384 wl_1_55
* net 385 wl_0_63
* net 390 rbl_wl_1_1
* net 391 wl_1_63
* net 392 wl_1_62
* net 393 vdd
* net 394 gnd
* cell instance $3 r0 *1 0,1.745
X$3 3 11 5 10 4 9 7 12 1 16 2 15 8 14 6 13 36 41 33 39 31 45 32 40 34 42 35 44
+ 37 43 38 71 66 68 63 75 62 74 64 69 65 70 61 73 67 72 96 101 94 102 92 103 98
+ 105 97 99 91 104 93 106 95 100 121 124 122 123 271 278 272 282 277 281 276
+ 280 275 285 265 291 266 290 268 288 270 286 269 287 267 289 264 292 263 279
+ 274 283 273 284 326 331 327 338 324 334 330 335 329 336 325 332 328 333 323
+ 337 356 362 361 363 359 368 357 367 354 366 355 365 358 364 360 387 385 386
+ 393 394 custom_sram_1r1w_32_256_freepdk45_wordline_buffer_array
* cell instance $18 r0 *1 6.3325,0
X$18 52 102 11 75 74 76 107 45 69 108 81 103 70 73 46 49 71 50 43 44 48 82 68
+ 79 101 42 40 72 53 78 77 80 112 39 19 10 9 21 22 12 16 23 20 15 14 51 47 41
+ 13 17 18 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179
+ 180 181 182 183 184 185 186 187 188 189 190 258 257 124 123 100 106 110 109
+ 104 105 99 259 111 113 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 331 340 388 345
+ 376 343 284 363 297 332 283 334 333 282 339 335 346 342 336 341 344 337 365
+ 305 338 362 372 281 370 374 369 298 366 306 387 285 295 296 287 278 371 286
+ 307 367 304 288 291 300 290 301 302 364 375 289 279 294 280 293 389 292 299
+ 373 368 386 303 393 394
+ custom_sram_1r1w_32_256_freepdk45_capped_replica_bitcell_array
* cell instance $19 r180 *1 55.66,100.415
X$19 390 388 391 389 392 371 380 373 381 370 379 369 382 375 383 374 378 376
+ 384 372 377 342 347 339 352 340 350 345 349 346 351 341 353 343 348 344 309
+ 297 313 296 308 294 322 293 314 298 318 295 319 307 316 304 315 301 321 300
+ 320 306 312 303 310 305 311 299 317 302 262 258 261 257 260 259 117 110 116
+ 109 119 111 118 113 114 108 120 107 115 112 85 78 90 77 87 76 86 82 88 81 89
+ 80 83 79 84 49 55 50 60 48 59 46 58 53 57 52 56 51 54 47 26 17 30 18 28 20 29
+ 23 27 22 24 21 25 19 393 394
+ custom_sram_1r1w_32_256_freepdk45_wordline_buffer_array
.ENDS custom_sram_1r1w_32_256_freepdk45_local_bitcell_array

* cell custom_sram_1r1w_32_256_freepdk45_pinv_16
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_16 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.275 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=3.6U AS=0.4095P AD=0.4095P PS=6.63U PD=6.63U
* device instance $13 r0 *1 0.2325,1.895 PMOS_VTG
M$13 3 1 2 3 PMOS_VTG L=0.05U W=10.8U AS=1.2285P AD=1.2285P PS=14.43U PD=14.43U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_16

* cell custom_sram_1r1w_32_256_freepdk45_pinv_17
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_17 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.2685 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=2.875U AS=0.32775P AD=0.32775P PS=5.4425U
+ PD=5.4425U
* device instance $11 r0 *1 0.2325,1.9125 PMOS_VTG
M$11 3 1 2 3 PMOS_VTG L=0.05U W=8.65U AS=0.9861P AD=0.9861P PS=11.795U
+ PD=11.795U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_17

* cell custom_sram_1r1w_32_256_freepdk45_pinv_7
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_7 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.26 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=1.08U AS=0.12555P AD=0.12555P PS=2.28U PD=2.28U
* device instance $5 r0 *1 0.2325,1.94 PMOS_VTG
M$5 3 1 2 3 PMOS_VTG L=0.05U W=3.24U AS=0.37665P AD=0.37665P PS=4.98U PD=4.98U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_7

* cell custom_sram_1r1w_32_256_freepdk45_pinv_6
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_6 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.215 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.36U AS=0.0432P AD=0.0432P PS=1.02U PD=1.02U
* device instance $3 r0 *1 0.2325,2.075 PMOS_VTG
M$3 3 1 2 3 PMOS_VTG L=0.05U W=1.08U AS=0.1296P AD=0.1296P PS=2.1U PD=2.1U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_6

* cell custom_sram_1r1w_32_256_freepdk45_pinv_5
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_5 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.215 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.02295P PS=0.615U PD=0.615U
* device instance $2 r0 *1 0.2325,2.075 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.54U AS=0.06885P AD=0.06885P PS=1.335U PD=1.335U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_5

* cell dff
* pin Q
* pin D
* pin clk
* pin vdd
* pin gnd
.SUBCKT dff 2 5 7 16 17
* net 2 Q
* net 5 D
* net 7 clk
* net 16 vdd
* net 17 gnd
* device instance $1 r0 *1 0.2925,1.5425 PMOS_VTG
M$1 16 5 13 16 PMOS_VTG L=0.05U W=0.5U AS=0.0525P AD=0.035P PS=1.21U PD=0.64U
* device instance $2 r0 *1 0.4825,1.5425 PMOS_VTG
M$2 13 7 4 16 PMOS_VTG L=0.05U W=0.5U AS=0.035P AD=0.035P PS=0.64U PD=0.64U
* device instance $3 r0 *1 0.6725,1.5425 PMOS_VTG
M$3 4 1 14 16 PMOS_VTG L=0.05U W=0.5U AS=0.035P AD=0.035P PS=0.64U PD=0.64U
* device instance $4 r0 *1 0.8625,1.5425 PMOS_VTG
M$4 14 6 16 16 PMOS_VTG L=0.05U W=0.5U AS=0.035P AD=0.0851P PS=0.64U PD=1.275U
* device instance $5 r0 *1 1.1575,1.5425 PMOS_VTG
M$5 16 4 6 16 PMOS_VTG L=0.05U W=0.5U AS=0.0851P AD=0.0525P PS=1.275U PD=1.21U
* device instance $6 r0 *1 2.2325,1.4525 PMOS_VTG
M$6 8 7 12 16 PMOS_VTG L=0.05U W=0.25U AS=0.038125P AD=0.0375P PS=0.7U PD=0.8U
* device instance $7 r0 *1 1.7925,1.5775 PMOS_VTG
M$7 16 6 15 16 PMOS_VTG L=0.05U W=0.5U AS=0.0875P AD=0.035P PS=1.245U PD=0.64U
* device instance $8 r0 *1 1.9825,1.5775 PMOS_VTG
M$8 15 1 8 16 PMOS_VTG L=0.05U W=0.5U AS=0.035P AD=0.038125P PS=0.64U PD=0.7U
* device instance $9 r0 *1 1.4975,1.65 PMOS_VTG
M$9 1 7 16 16 PMOS_VTG L=0.05U W=1U AS=0.105P AD=0.0875P PS=2.21U PD=1.245U
* device instance $10 r0 *1 2.3225,2.0175 PMOS_VTG
M$10 16 2 12 16 PMOS_VTG L=0.05U W=0.25U AS=0.055125P AD=0.02625P PS=1.21U
+ PD=0.71U
* device instance $11 r0 *1 2.5825,1.7925 PMOS_VTG
M$11 16 8 2 16 PMOS_VTG L=0.05U W=1U AS=0.055125P AD=0.105P PS=1.21U PD=2.21U
* device instance $12 r0 *1 2.0475,0.3475 NMOS_VTG
M$12 17 2 3 17 NMOS_VTG L=0.05U W=0.25U AS=0.02625P AD=0.02625P PS=0.71U
+ PD=0.71U
* device instance $13 r0 *1 2.5825,0.7125 NMOS_VTG
M$13 17 8 2 17 NMOS_VTG L=0.05U W=0.5U AS=0.0775P AD=0.0525P PS=1.31U PD=1.21U
* device instance $14 r0 *1 0.2925,0.725 NMOS_VTG
M$14 17 5 9 17 NMOS_VTG L=0.05U W=0.25U AS=0.02625P AD=0.0175P PS=0.71U PD=0.39U
* device instance $15 r0 *1 0.4825,0.725 NMOS_VTG
M$15 9 1 4 17 NMOS_VTG L=0.05U W=0.25U AS=0.0175P AD=0.0175P PS=0.39U PD=0.39U
* device instance $16 r0 *1 0.6725,0.725 NMOS_VTG
M$16 4 7 10 17 NMOS_VTG L=0.05U W=0.25U AS=0.0175P AD=0.0175P PS=0.39U PD=0.39U
* device instance $17 r0 *1 0.8625,0.725 NMOS_VTG
M$17 17 6 10 17 NMOS_VTG L=0.05U W=0.25U AS=0.0502P AD=0.0175P PS=0.93U PD=0.39U
* device instance $18 r0 *1 1.1575,0.725 NMOS_VTG
M$18 17 4 6 17 NMOS_VTG L=0.05U W=0.25U AS=0.0502P AD=0.02625P PS=0.93U PD=0.71U
* device instance $19 r0 *1 1.4975,0.6575 NMOS_VTG
M$19 1 7 17 17 NMOS_VTG L=0.05U W=0.5U AS=0.0525P AD=0.04375P PS=1.21U PD=0.745U
* device instance $20 r0 *1 1.7925,0.7825 NMOS_VTG
M$20 17 6 11 17 NMOS_VTG L=0.05U W=0.25U AS=0.04375P AD=0.0175P PS=0.745U
+ PD=0.39U
* device instance $21 r0 *1 1.9825,0.7825 NMOS_VTG
M$21 11 7 8 17 NMOS_VTG L=0.05U W=0.25U AS=0.0175P AD=0.0175P PS=0.39U PD=0.39U
* device instance $22 r0 *1 2.1725,0.7825 NMOS_VTG
M$22 8 1 3 17 NMOS_VTG L=0.05U W=0.25U AS=0.0175P AD=0.0275P PS=0.39U PD=0.72U
.ENDS dff

* cell custom_sram_1r1w_32_256_freepdk45_pand2
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pand2 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0,0
X$1 3 4 1 5 6 custom_sram_1r1w_32_256_freepdk45_pnand2_0
* cell instance $2 r0 *1 0.75,0
X$2 2 1 5 6 custom_sram_1r1w_32_256_freepdk45_pdriver
.ENDS custom_sram_1r1w_32_256_freepdk45_pand2

* cell custom_sram_1r1w_32_256_freepdk45_pinv_4
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_4 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.17 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.09U AS=0.011475P AD=0.011475P PS=0.435U
+ PD=0.435U
* device instance $2 r0 *1 0.2325,2.21 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_4

* cell custom_sram_1r1w_32_256_freepdk45_wordline_driver
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_wordline_driver 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0.9025,0
X$1 2 1 5 6 custom_sram_1r1w_32_256_freepdk45_pbuf
* cell instance $2 r0 *1 0,0
X$2 3 4 1 5 6 custom_sram_1r1w_32_256_freepdk45_pnand2
.ENDS custom_sram_1r1w_32_256_freepdk45_wordline_driver

* cell custom_sram_1r1w_32_256_freepdk45_hierarchical_predecode2x4
* pin in_0
* pin in_1
* pin out_0
* pin out_1
* pin out_2
* pin out_3
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_hierarchical_predecode2x4 1 2 5 6 7 8
+ 9 10
* net 1 in_0
* net 2 in_1
* net 5 out_0
* net 6 out_1
* net 7 out_2
* net 8 out_3
* net 9 vdd
* net 10 gnd
* cell instance $1 m0 *1 2.0875,2.99
X$1 6 1 4 9 10 custom_sram_1r1w_32_256_freepdk45_and2_dec
* cell instance $2 m0 *1 2.0875,5.98
X$2 8 1 2 9 10 custom_sram_1r1w_32_256_freepdk45_and2_dec
* cell instance $8 r0 *1 0.56,0
X$8 1 3 9 10 custom_sram_1r1w_32_256_freepdk45_pinv_0
* cell instance $9 r0 *1 2.0875,2.99
X$9 7 3 2 9 10 custom_sram_1r1w_32_256_freepdk45_and2_dec
* cell instance $15 m0 *1 0.56,2.99
X$15 2 4 9 10 custom_sram_1r1w_32_256_freepdk45_pinv_0
* cell instance $16 r0 *1 2.0875,0
X$16 5 3 4 9 10 custom_sram_1r1w_32_256_freepdk45_and2_dec
.ENDS custom_sram_1r1w_32_256_freepdk45_hierarchical_predecode2x4

* cell custom_sram_1r1w_32_256_freepdk45_and3_dec
* pin Z
* pin A
* pin B
* pin C
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_and3_dec 2 3 4 5 6 7
* net 2 Z
* net 3 A
* net 4 B
* net 5 C
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 0,0
X$1 3 4 5 1 6 7 custom_sram_1r1w_32_256_freepdk45_pnand3
* cell instance $2 r0 *1 1.2475,0
X$2 1 2 6 7 custom_sram_1r1w_32_256_freepdk45_pinv_0
.ENDS custom_sram_1r1w_32_256_freepdk45_and3_dec

* cell custom_sram_1r1w_32_256_freepdk45_column_mux_0
* pin sel
* pin bl
* pin br_out
* pin bl_out
* pin br
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_column_mux_0 1 2 3 4 5 6
* net 1 sel
* net 2 bl
* net 3 br_out
* net 4 bl_out
* net 5 br
* net 6 gnd
* device instance $1 r0 *1 0.5875,0.44 NMOS_VTG
M$1 3 1 5 6 NMOS_VTG L=0.05U W=0.72U AS=0.0918P AD=0.0918P PS=1.695U PD=1.695U
* device instance $2 r0 *1 0.5875,1.3 NMOS_VTG
M$2 4 1 2 6 NMOS_VTG L=0.05U W=0.72U AS=0.0918P AD=0.0918P PS=1.695U PD=1.695U
.ENDS custom_sram_1r1w_32_256_freepdk45_column_mux_0

* cell sense_amp
* pin br
* pin dout
* pin bl
* pin en
* pin vdd
* pin gnd
.SUBCKT sense_amp 1 3 4 6 9 10
* net 1 br
* net 3 dout
* net 4 bl
* net 6 en
* net 9 vdd
* net 10 gnd
* device instance $1 r0 *1 0.2575,4.0975 PMOS_VTG
M$1 5 7 9 9 PMOS_VTG L=0.05U W=0.54U AS=0.0567P AD=0.0378P PS=1.29U PD=0.68U
* device instance $2 r0 *1 0.4475,4.0975 PMOS_VTG
M$2 9 5 7 9 PMOS_VTG L=0.05U W=0.54U AS=0.0378P AD=0.0567P PS=0.68U PD=1.29U
* device instance $3 r0 *1 0.4475,3.15 PMOS_VTG
M$3 7 6 1 9 PMOS_VTG L=0.05U W=0.72U AS=0.0756P AD=0.0756P PS=1.65U PD=1.65U
* device instance $4 r0 *1 0.2575,2.18 PMOS_VTG
M$4 4 6 5 9 PMOS_VTG L=0.05U W=0.72U AS=0.0756P AD=0.0756P PS=1.65U PD=1.65U
* device instance $5 r0 *1 0.4625,0.955 PMOS_VTG
M$5 9 5 2 9 PMOS_VTG L=0.05U W=0.18U AS=0.03285P AD=0.0189P PS=0.695U PD=0.57U
* device instance $6 r0 *1 0.2575,1.135 PMOS_VTG
M$6 3 2 9 9 PMOS_VTG L=0.05U W=0.54U AS=0.0567P AD=0.03285P PS=1.29U PD=0.695U
* device instance $7 r0 *1 0.3575,5.445 NMOS_VTG
M$7 8 6 10 10 NMOS_VTG L=0.05U W=0.27U AS=0.02835P AD=0.02835P PS=0.75U PD=0.75U
* device instance $8 r0 *1 0.2575,4.9875 NMOS_VTG
M$8 5 7 8 10 NMOS_VTG L=0.05U W=0.27U AS=0.02835P AD=0.0189P PS=0.75U PD=0.41U
* device instance $9 r0 *1 0.4475,4.9875 NMOS_VTG
M$9 8 5 7 10 NMOS_VTG L=0.05U W=0.27U AS=0.0189P AD=0.02835P PS=0.41U PD=0.75U
* device instance $10 r0 *1 0.2575,0.245 NMOS_VTG
M$10 3 2 10 10 NMOS_VTG L=0.05U W=0.27U AS=0.02835P AD=0.016425P PS=0.75U
+ PD=0.425U
* device instance $11 r0 *1 0.4625,0.335 NMOS_VTG
M$11 10 5 2 10 NMOS_VTG L=0.05U W=0.09U AS=0.016425P AD=0.00945P PS=0.425U
+ PD=0.39U
.ENDS sense_amp

* cell custom_sram_1r1w_32_256_freepdk45_precharge_1
* pin en_bar
* pin bl
* pin br
* pin vdd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_precharge_1 1 2 3 4
* net 1 en_bar
* net 2 bl
* net 3 br
* net 4 vdd
* device instance $1 r0 *1 0.265,0.905 PMOS_VTG
M$1 2 1 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.48,0.905 PMOS_VTG
M$2 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.265,0.355 PMOS_VTG
M$3 2 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS custom_sram_1r1w_32_256_freepdk45_precharge_1

* cell custom_sram_1r1w_32_256_freepdk45_column_mux
* pin sel
* pin bl
* pin br_out
* pin bl_out
* pin br
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_column_mux 1 2 3 4 5 6
* net 1 sel
* net 2 bl
* net 3 br_out
* net 4 bl_out
* net 5 br
* net 6 gnd
* device instance $1 r0 *1 0.5875,1.3 NMOS_VTG
M$1 4 1 2 6 NMOS_VTG L=0.05U W=0.72U AS=0.0918P AD=0.0918P PS=1.695U PD=1.695U
* device instance $2 r0 *1 0.5875,0.44 NMOS_VTG
M$2 3 1 5 6 NMOS_VTG L=0.05U W=0.72U AS=0.0918P AD=0.0918P PS=1.695U PD=1.695U
.ENDS custom_sram_1r1w_32_256_freepdk45_column_mux

* cell write_driver
* pin din
* pin en
* pin br
* pin bl
* pin vdd
* pin gnd
.SUBCKT write_driver 1 2 5 9 11 12
* net 1 din
* net 2 en
* net 5 br
* net 9 bl
* net 11 vdd
* net 12 gnd
* device instance $1 r0 *1 0.17,3.0725 PMOS_VTG
M$1 11 3 8 11 PMOS_VTG L=0.05U W=0.36U AS=0.0378P AD=0.0252P PS=0.93U PD=0.5U
* device instance $2 r0 *1 0.36,3.0725 PMOS_VTG
M$2 8 4 9 11 PMOS_VTG L=0.05U W=0.36U AS=0.0252P AD=0.0378P PS=0.5U PD=0.93U
* device instance $3 r0 *1 0.17,2.46 PMOS_VTG
M$3 11 1 7 11 PMOS_VTG L=0.05U W=0.36U AS=0.0378P AD=0.0252P PS=0.93U PD=0.5U
* device instance $4 r0 *1 0.36,2.46 PMOS_VTG
M$4 7 4 5 11 PMOS_VTG L=0.05U W=0.36U AS=0.0252P AD=0.0378P PS=0.5U PD=0.93U
* device instance $5 r0 *1 0.51,0.885 PMOS_VTG
M$5 4 2 11 11 PMOS_VTG L=0.05U W=0.36U AS=0.0378P AD=0.0378P PS=0.93U PD=0.93U
* device instance $6 r0 *1 0.17,0.885 PMOS_VTG
M$6 11 1 3 11 PMOS_VTG L=0.05U W=0.36U AS=0.0378P AD=0.0378P PS=0.93U PD=0.93U
* device instance $7 r0 *1 0.17,3.6775 NMOS_VTG
M$7 12 3 10 12 NMOS_VTG L=0.05U W=0.18U AS=0.0189P AD=0.0126P PS=0.57U PD=0.32U
* device instance $8 r0 *1 0.36,3.6775 NMOS_VTG
M$8 10 2 9 12 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.0189P PS=0.32U PD=0.57U
* device instance $9 r0 *1 0.17,1.855 NMOS_VTG
M$9 12 1 6 12 NMOS_VTG L=0.05U W=0.18U AS=0.0189P AD=0.0126P PS=0.57U PD=0.32U
* device instance $10 r0 *1 0.36,1.855 NMOS_VTG
M$10 6 2 5 12 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.0189P PS=0.32U PD=0.57U
* device instance $11 r0 *1 0.51,1.49 NMOS_VTG
M$11 4 2 12 12 NMOS_VTG L=0.05U W=0.18U AS=0.0189P AD=0.0189P PS=0.57U PD=0.57U
* device instance $12 r0 *1 0.17,1.49 NMOS_VTG
M$12 12 1 3 12 NMOS_VTG L=0.05U W=0.18U AS=0.0189P AD=0.0189P PS=0.57U PD=0.57U
.ENDS write_driver

* cell custom_sram_1r1w_32_256_freepdk45_precharge_0
* pin en_bar
* pin bl
* pin br
* pin vdd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_precharge_0 1 2 3 4
* net 1 en_bar
* net 2 bl
* net 3 br
* net 4 vdd
* device instance $1 r0 *1 0.265,0.905 PMOS_VTG
M$1 2 1 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.48,0.905 PMOS_VTG
M$2 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.265,0.355 PMOS_VTG
M$3 2 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS custom_sram_1r1w_32_256_freepdk45_precharge_0

* cell custom_sram_1r1w_32_256_freepdk45_capped_replica_bitcell_array_1
* pin wl_1_9
* pin wl_0_23
* pin rbl_wl_0_0
* pin wl_0_16
* pin wl_0_17
* pin wl_1_19
* pin wl_1_23
* pin wl_0_9
* pin wl_0_18
* pin wl_1_24
* pin wl_1_17
* pin wl_0_24
* pin wl_0_19
* pin wl_0_20
* pin wl_1_11
* pin wl_1_14
* pin wl_0_14
* pin wl_1_13
* pin wl_0_13
* pin wl_0_12
* pin wl_1_12
* pin wl_1_18
* pin wl_0_15
* pin wl_1_15
* pin wl_0_22
* pin wl_0_11
* pin wl_0_10
* pin wl_0_21
* pin wl_1_10
* pin wl_1_21
* pin wl_1_20
* pin wl_1_16
* pin wl_1_22
* pin wl_0_8
* pin wl_1_0
* pin wl_0_0
* pin wl_0_1
* pin wl_1_1
* pin wl_1_2
* pin wl_0_2
* pin wl_0_3
* pin wl_1_3
* pin wl_1_4
* pin wl_0_4
* pin wl_0_5
* pin wl_1_8
* pin wl_1_7
* pin wl_0_7
* pin wl_0_6
* pin wl_1_6
* pin wl_1_5
* pin bl_0_0
* pin bl_1_0
* pin br_1_0
* pin br_0_0
* pin bl_0_1
* pin bl_1_1
* pin br_1_1
* pin br_0_1
* pin bl_0_2
* pin bl_1_2
* pin br_1_2
* pin br_0_2
* pin bl_0_3
* pin bl_1_3
* pin br_1_3
* pin br_0_3
* pin bl_0_4
* pin bl_1_4
* pin br_1_4
* pin br_0_4
* pin bl_0_5
* pin bl_1_5
* pin br_1_5
* pin br_0_5
* pin bl_0_6
* pin bl_1_6
* pin br_1_6
* pin br_0_6
* pin bl_0_7
* pin bl_1_7
* pin br_1_7
* pin br_0_7
* pin bl_0_8
* pin bl_1_8
* pin br_1_8
* pin br_0_8
* pin bl_0_9
* pin bl_1_9
* pin br_1_9
* pin br_0_9
* pin bl_0_10
* pin bl_1_10
* pin br_1_10
* pin br_0_10
* pin bl_0_11
* pin bl_1_11
* pin br_1_11
* pin br_0_11
* pin bl_0_12
* pin bl_1_12
* pin br_1_12
* pin br_0_12
* pin bl_0_13
* pin bl_1_13
* pin br_1_13
* pin br_0_13
* pin bl_0_14
* pin bl_1_14
* pin br_1_14
* pin br_0_14
* pin bl_0_15
* pin bl_1_15
* pin br_1_15
* pin br_0_15
* pin bl_0_16
* pin bl_1_16
* pin wl_1_31
* pin wl_1_30
* pin wl_0_30
* pin wl_0_31
* pin wl_0_29
* pin wl_0_28
* pin wl_1_28
* pin wl_1_27
* pin wl_0_27
* pin wl_0_25
* pin wl_0_26
* pin wl_1_29
* pin wl_1_26
* pin wl_1_25
* pin br_1_16
* pin br_0_16
* pin bl_0_17
* pin bl_1_17
* pin br_1_17
* pin br_0_17
* pin bl_0_18
* pin bl_1_18
* pin br_1_18
* pin br_0_18
* pin bl_0_19
* pin bl_1_19
* pin br_1_19
* pin br_0_19
* pin bl_0_20
* pin bl_1_20
* pin br_1_20
* pin br_0_20
* pin bl_0_21
* pin bl_1_21
* pin br_1_21
* pin br_0_21
* pin bl_0_22
* pin bl_1_22
* pin br_1_22
* pin br_0_22
* pin bl_0_23
* pin bl_1_23
* pin br_1_23
* pin br_0_23
* pin bl_0_24
* pin bl_1_24
* pin br_1_24
* pin br_0_24
* pin bl_0_25
* pin bl_1_25
* pin br_1_25
* pin br_0_25
* pin bl_0_26
* pin bl_1_26
* pin br_1_26
* pin br_0_26
* pin bl_0_27
* pin bl_1_27
* pin br_1_27
* pin br_0_27
* pin bl_0_28
* pin bl_1_28
* pin br_1_28
* pin br_0_28
* pin bl_0_29
* pin bl_1_29
* pin br_1_29
* pin br_0_29
* pin bl_0_30
* pin bl_1_30
* pin br_1_30
* pin br_0_30
* pin bl_0_31
* pin bl_1_31
* pin br_1_31
* pin br_0_31
* pin rbl_bl_0_1
* pin rbl_bl_1_1
* pin rbl_br_1_1
* pin rbl_br_0_1
* pin wl_0_47
* pin wl_1_52
* pin rbl_wl_1_1
* pin wl_1_51
* pin wl_1_56
* pin wl_1_48
* pin wl_0_46
* pin wl_0_56
* pin wl_1_46
* pin wl_0_52
* pin wl_0_45
* pin wl_0_49
* pin wl_0_53
* pin wl_0_33
* pin wl_1_53
* pin wl_0_50
* pin wl_1_50
* pin wl_1_54
* pin wl_0_51
* pin wl_1_49
* pin wl_1_47
* pin wl_0_54
* pin wl_0_60
* pin wl_1_34
* pin wl_0_48
* pin wl_0_55
* pin wl_1_55
* pin wl_0_34
* pin wl_1_60
* pin wl_1_57
* pin wl_1_59
* pin wl_1_42
* pin wl_0_59
* pin wl_1_36
* pin wl_0_62
* pin wl_0_36
* pin wl_1_41
* pin wl_1_45
* pin wl_0_41
* pin wl_0_32
* pin wl_1_62
* pin wl_0_40
* pin wl_1_40
* pin wl_0_58
* pin wl_1_39
* pin wl_0_39
* pin wl_0_37
* pin wl_1_37
* pin wl_0_38
* pin wl_1_38
* pin wl_1_32
* pin wl_0_61
* pin wl_1_58
* pin wl_0_42
* pin wl_0_44
* pin wl_1_44
* pin wl_0_35
* pin wl_1_43
* pin wl_1_63
* pin wl_0_43
* pin wl_1_33
* pin wl_1_61
* pin wl_0_57
* pin wl_0_63
* pin wl_1_35
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_capped_replica_bitcell_array_1 1 2 3
+ 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31
+ 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57
+ 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106
+ 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125
+ 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144
+ 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239
+ 240 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258
+ 259 260 261 262 263 264
* net 1 wl_1_9
* net 2 wl_0_23
* net 3 rbl_wl_0_0
* net 4 wl_0_16
* net 5 wl_0_17
* net 6 wl_1_19
* net 7 wl_1_23
* net 8 wl_0_9
* net 9 wl_0_18
* net 10 wl_1_24
* net 11 wl_1_17
* net 12 wl_0_24
* net 13 wl_0_19
* net 14 wl_0_20
* net 15 wl_1_11
* net 16 wl_1_14
* net 17 wl_0_14
* net 18 wl_1_13
* net 19 wl_0_13
* net 20 wl_0_12
* net 21 wl_1_12
* net 22 wl_1_18
* net 23 wl_0_15
* net 24 wl_1_15
* net 25 wl_0_22
* net 26 wl_0_11
* net 27 wl_0_10
* net 28 wl_0_21
* net 29 wl_1_10
* net 30 wl_1_21
* net 31 wl_1_20
* net 32 wl_1_16
* net 33 wl_1_22
* net 34 wl_0_8
* net 35 wl_1_0
* net 36 wl_0_0
* net 37 wl_0_1
* net 38 wl_1_1
* net 39 wl_1_2
* net 40 wl_0_2
* net 41 wl_0_3
* net 42 wl_1_3
* net 43 wl_1_4
* net 44 wl_0_4
* net 45 wl_0_5
* net 46 wl_1_8
* net 47 wl_1_7
* net 48 wl_0_7
* net 49 wl_0_6
* net 50 wl_1_6
* net 51 wl_1_5
* net 52 bl_0_0
* net 53 bl_1_0
* net 54 br_1_0
* net 55 br_0_0
* net 56 bl_0_1
* net 57 bl_1_1
* net 58 br_1_1
* net 59 br_0_1
* net 60 bl_0_2
* net 61 bl_1_2
* net 62 br_1_2
* net 63 br_0_2
* net 64 bl_0_3
* net 65 bl_1_3
* net 66 br_1_3
* net 67 br_0_3
* net 68 bl_0_4
* net 69 bl_1_4
* net 70 br_1_4
* net 71 br_0_4
* net 72 bl_0_5
* net 73 bl_1_5
* net 74 br_1_5
* net 75 br_0_5
* net 76 bl_0_6
* net 77 bl_1_6
* net 78 br_1_6
* net 79 br_0_6
* net 80 bl_0_7
* net 81 bl_1_7
* net 82 br_1_7
* net 83 br_0_7
* net 84 bl_0_8
* net 85 bl_1_8
* net 86 br_1_8
* net 87 br_0_8
* net 88 bl_0_9
* net 89 bl_1_9
* net 90 br_1_9
* net 91 br_0_9
* net 92 bl_0_10
* net 93 bl_1_10
* net 94 br_1_10
* net 95 br_0_10
* net 96 bl_0_11
* net 97 bl_1_11
* net 98 br_1_11
* net 99 br_0_11
* net 100 bl_0_12
* net 101 bl_1_12
* net 102 br_1_12
* net 103 br_0_12
* net 104 bl_0_13
* net 105 bl_1_13
* net 106 br_1_13
* net 107 br_0_13
* net 108 bl_0_14
* net 109 bl_1_14
* net 110 br_1_14
* net 111 br_0_14
* net 112 bl_0_15
* net 113 bl_1_15
* net 114 br_1_15
* net 115 br_0_15
* net 116 bl_0_16
* net 117 bl_1_16
* net 118 wl_1_31
* net 119 wl_1_30
* net 120 wl_0_30
* net 121 wl_0_31
* net 122 wl_0_29
* net 123 wl_0_28
* net 124 wl_1_28
* net 125 wl_1_27
* net 126 wl_0_27
* net 127 wl_0_25
* net 128 wl_0_26
* net 129 wl_1_29
* net 130 wl_1_26
* net 131 wl_1_25
* net 132 br_1_16
* net 133 br_0_16
* net 134 bl_0_17
* net 135 bl_1_17
* net 136 br_1_17
* net 137 br_0_17
* net 138 bl_0_18
* net 139 bl_1_18
* net 140 br_1_18
* net 141 br_0_18
* net 142 bl_0_19
* net 143 bl_1_19
* net 144 br_1_19
* net 145 br_0_19
* net 146 bl_0_20
* net 147 bl_1_20
* net 148 br_1_20
* net 149 br_0_20
* net 150 bl_0_21
* net 151 bl_1_21
* net 152 br_1_21
* net 153 br_0_21
* net 154 bl_0_22
* net 155 bl_1_22
* net 156 br_1_22
* net 157 br_0_22
* net 158 bl_0_23
* net 159 bl_1_23
* net 160 br_1_23
* net 161 br_0_23
* net 162 bl_0_24
* net 163 bl_1_24
* net 164 br_1_24
* net 165 br_0_24
* net 166 bl_0_25
* net 167 bl_1_25
* net 168 br_1_25
* net 169 br_0_25
* net 170 bl_0_26
* net 171 bl_1_26
* net 172 br_1_26
* net 173 br_0_26
* net 174 bl_0_27
* net 175 bl_1_27
* net 176 br_1_27
* net 177 br_0_27
* net 178 bl_0_28
* net 179 bl_1_28
* net 180 br_1_28
* net 181 br_0_28
* net 182 bl_0_29
* net 183 bl_1_29
* net 184 br_1_29
* net 185 br_0_29
* net 186 bl_0_30
* net 187 bl_1_30
* net 188 br_1_30
* net 189 br_0_30
* net 190 bl_0_31
* net 191 bl_1_31
* net 192 br_1_31
* net 193 br_0_31
* net 194 rbl_bl_0_1
* net 195 rbl_bl_1_1
* net 196 rbl_br_1_1
* net 197 rbl_br_0_1
* net 198 wl_0_47
* net 199 wl_1_52
* net 200 rbl_wl_1_1
* net 201 wl_1_51
* net 202 wl_1_56
* net 203 wl_1_48
* net 204 wl_0_46
* net 205 wl_0_56
* net 206 wl_1_46
* net 207 wl_0_52
* net 208 wl_0_45
* net 209 wl_0_49
* net 210 wl_0_53
* net 211 wl_0_33
* net 212 wl_1_53
* net 213 wl_0_50
* net 214 wl_1_50
* net 215 wl_1_54
* net 216 wl_0_51
* net 217 wl_1_49
* net 218 wl_1_47
* net 219 wl_0_54
* net 220 wl_0_60
* net 221 wl_1_34
* net 222 wl_0_48
* net 223 wl_0_55
* net 224 wl_1_55
* net 225 wl_0_34
* net 226 wl_1_60
* net 227 wl_1_57
* net 228 wl_1_59
* net 229 wl_1_42
* net 230 wl_0_59
* net 231 wl_1_36
* net 232 wl_0_62
* net 233 wl_0_36
* net 234 wl_1_41
* net 235 wl_1_45
* net 236 wl_0_41
* net 237 wl_0_32
* net 238 wl_1_62
* net 239 wl_0_40
* net 240 wl_1_40
* net 241 wl_0_58
* net 242 wl_1_39
* net 243 wl_0_39
* net 244 wl_0_37
* net 245 wl_1_37
* net 246 wl_0_38
* net 247 wl_1_38
* net 248 wl_1_32
* net 249 wl_0_61
* net 250 wl_1_58
* net 251 wl_0_42
* net 252 wl_0_44
* net 253 wl_1_44
* net 254 wl_0_35
* net 255 wl_1_43
* net 256 wl_1_63
* net 257 wl_0_43
* net 258 wl_1_33
* net 259 wl_1_61
* net 260 wl_0_57
* net 261 wl_0_63
* net 262 wl_1_35
* net 263 vdd
* net 264 gnd
* cell instance $1 r0 *1 2.11,1.745
X$1 264 3 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74
+ 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99
+ 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 132
+ 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151
+ 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170
+ 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189
+ 190 191 192 193 194 195 196 197 36 35 38 37 39 40 42 41 43 44 51 45 49 50 47
+ 48 34 46 1 8 29 27 15 26 21 20 18 19 17 16 24 23 4 32 11 5 9 22 6 13 14 31 30
+ 28 25 33 7 2 12 10 131 127 128 130 125 126 123 124 129 122 120 119 118 121
+ 237 248 211 258 225 221 262 254 233 231 245 244 246 247 242 243 239 240 236
+ 234 251 229 257 255 253 252 208 235 204 206 218 198 222 203 217 209 213 214
+ 216 201 207 199 210 212 215 219 224 223 205 202 227 260 241 250 228 230 220
+ 226 259 249 232 238 256 261 264 200 263 264
+ custom_sram_1r1w_32_256_freepdk45_replica_bitcell_array_1
* cell instance $2 r0 *1 0.935,0.25
X$2 264 264 3 264 35 36 37 38 39 40 41 42 43 44 45 51 50 49 48 47 46 34 8 1 29
+ 27 26 15 21 20 19 18 16 17 23 24 32 4 5 11 22 9 13 6 31 14 28 30 33 25 2 7 10
+ 12 127 131 130 128 126 125 124 123 122 129 119 120 121 118 248 237 211 258
+ 221 225 254 262 231 233 244 245 247 246 243 242 240 239 236 234 229 251 257
+ 255 253 252 208 235 206 204 198 218 203 222 209 217 214 213 216 201 199 207
+ 210 212 215 219 223 224 202 205 260 227 250 241 230 228 226 220 249 259 238
+ 232 261 256 200 264 264 264 263 264
+ custom_sram_1r1w_32_256_freepdk45_dummy_array_2
* cell instance $3 r0 *1 40.885,0.25
X$3 264 264 3 264 35 36 37 38 39 40 41 42 43 44 45 51 50 49 48 47 46 34 8 1 29
+ 27 26 15 21 20 19 18 16 17 23 24 32 4 5 11 22 9 13 6 31 14 28 30 33 25 2 7 10
+ 12 127 131 130 128 126 125 124 123 122 129 119 120 121 118 248 237 211 258
+ 221 225 254 262 231 233 244 245 247 246 243 242 240 239 236 234 229 251 257
+ 255 253 252 208 235 206 204 198 218 203 222 209 217 214 213 216 201 199 207
+ 210 212 215 219 223 224 202 205 260 227 250 241 230 228 226 220 249 259 238
+ 232 261 256 200 264 264 264 263 264
+ custom_sram_1r1w_32_256_freepdk45_dummy_array_7
* cell instance $4 r0 *1 2.11,0.25
X$4 264 264 263 264 custom_sram_1r1w_32_256_freepdk45_dummy_array_1
* cell instance $5 m0 *1 2.11,101.91
X$5 264 264 263 264 custom_sram_1r1w_32_256_freepdk45_dummy_array_0
.ENDS custom_sram_1r1w_32_256_freepdk45_capped_replica_bitcell_array_1

* cell custom_sram_1r1w_32_256_freepdk45_capped_replica_bitcell_array_0
* pin wl_1_9
* pin wl_1_20
* pin wl_1_19
* pin wl_0_9
* pin wl_1_23
* pin wl_0_19
* pin wl_0_8
* pin wl_0_18
* pin wl_1_8
* pin wl_1_18
* pin wl_1_12
* pin wl_0_12
* pin wl_0_23
* pin wl_1_3
* pin wl_1_10
* pin wl_0_20
* pin wl_0_10
* pin wl_0_21
* pin wl_1_15
* pin wl_0_22
* pin wl_0_11
* pin wl_1_21
* pin wl_1_11
* pin wl_1_22
* pin wl_1_2
* pin wl_1_16
* pin wl_1_5
* pin wl_1_0
* pin wl_0_5
* pin wl_0_0
* pin wl_0_1
* pin wl_1_1
* pin wl_0_14
* pin wl_0_15
* pin wl_0_4
* pin wl_0_2
* pin wl_1_4
* pin wl_1_13
* pin wl_0_3
* pin wl_0_13
* pin wl_0_16
* pin wl_1_7
* pin wl_1_14
* pin wl_0_7
* pin wl_1_6
* pin rbl_wl_0_0
* pin wl_0_6
* pin wl_0_17
* pin wl_1_17
* pin bl_0_0
* pin bl_1_0
* pin br_1_0
* pin br_0_0
* pin bl_0_1
* pin bl_1_1
* pin br_1_1
* pin br_0_1
* pin bl_0_2
* pin bl_1_2
* pin br_1_2
* pin br_0_2
* pin bl_0_3
* pin bl_1_3
* pin br_1_3
* pin br_0_3
* pin bl_0_4
* pin bl_1_4
* pin br_1_4
* pin br_0_4
* pin bl_0_5
* pin bl_1_5
* pin br_1_5
* pin br_0_5
* pin bl_0_6
* pin bl_1_6
* pin br_1_6
* pin br_0_6
* pin bl_0_7
* pin bl_1_7
* pin br_1_7
* pin br_0_7
* pin bl_0_8
* pin bl_1_8
* pin br_1_8
* pin br_0_8
* pin bl_0_9
* pin bl_1_9
* pin br_1_9
* pin br_0_9
* pin bl_0_10
* pin bl_1_10
* pin br_1_10
* pin br_0_10
* pin bl_0_11
* pin bl_1_11
* pin br_1_11
* pin br_0_11
* pin bl_0_12
* pin bl_1_12
* pin br_1_12
* pin br_0_12
* pin bl_0_13
* pin bl_1_13
* pin br_1_13
* pin br_0_13
* pin bl_0_14
* pin bl_1_14
* pin br_1_14
* pin br_0_14
* pin bl_0_15
* pin bl_1_15
* pin br_1_15
* pin br_0_15
* pin wl_0_27
* pin wl_0_30
* pin wl_1_30
* pin wl_1_24
* pin wl_1_29
* pin wl_0_24
* pin wl_0_29
* pin wl_0_25
* pin wl_0_31
* pin wl_1_25
* pin wl_1_31
* pin wl_1_26
* pin wl_0_28
* pin wl_0_26
* pin wl_1_28
* pin wl_1_27
* pin bl_0_16
* pin bl_1_16
* pin br_1_16
* pin br_0_16
* pin bl_0_17
* pin bl_1_17
* pin br_1_17
* pin br_0_17
* pin bl_0_18
* pin bl_1_18
* pin br_1_18
* pin br_0_18
* pin bl_0_19
* pin bl_1_19
* pin br_1_19
* pin br_0_19
* pin bl_0_20
* pin bl_1_20
* pin br_1_20
* pin br_0_20
* pin bl_0_21
* pin bl_1_21
* pin br_1_21
* pin br_0_21
* pin bl_0_22
* pin bl_1_22
* pin br_1_22
* pin br_0_22
* pin bl_0_23
* pin bl_1_23
* pin br_1_23
* pin br_0_23
* pin bl_0_24
* pin bl_1_24
* pin br_1_24
* pin br_0_24
* pin bl_0_25
* pin bl_1_25
* pin br_1_25
* pin br_0_25
* pin bl_0_26
* pin bl_1_26
* pin br_1_26
* pin br_0_26
* pin bl_0_27
* pin bl_1_27
* pin br_1_27
* pin br_0_27
* pin bl_0_28
* pin bl_1_28
* pin br_1_28
* pin br_0_28
* pin bl_0_29
* pin bl_1_29
* pin br_1_29
* pin br_0_29
* pin bl_0_30
* pin bl_1_30
* pin br_1_30
* pin br_0_30
* pin bl_0_31
* pin bl_1_31
* pin br_1_31
* pin br_0_31
* pin wl_1_62
* pin wl_0_62
* pin rbl_wl_1_1
* pin wl_1_49
* pin wl_0_49
* pin wl_0_48
* pin wl_1_48
* pin wl_0_63
* pin wl_1_50
* pin wl_1_63
* pin wl_1_47
* pin wl_0_50
* pin wl_0_47
* pin wl_0_59
* pin wl_1_55
* pin wl_0_58
* pin wl_1_58
* pin wl_1_59
* pin wl_0_32
* pin wl_1_57
* pin wl_0_57
* pin wl_1_60
* pin wl_0_56
* pin wl_1_56
* pin wl_0_60
* pin wl_0_51
* pin wl_0_55
* pin wl_0_61
* pin wl_0_54
* pin wl_1_54
* pin wl_1_53
* pin wl_0_53
* pin wl_0_52
* pin wl_1_52
* pin wl_1_51
* pin wl_1_61
* pin wl_0_39
* pin wl_0_44
* pin wl_0_35
* pin wl_1_35
* pin wl_1_36
* pin wl_1_44
* pin wl_0_36
* pin wl_0_37
* pin wl_1_37
* pin wl_1_38
* pin wl_0_38
* pin wl_0_46
* pin wl_1_39
* pin wl_1_43
* pin wl_1_40
* pin wl_0_40
* pin wl_0_43
* pin wl_0_41
* pin wl_1_41
* pin wl_1_42
* pin wl_0_42
* pin wl_0_45
* pin wl_0_34
* pin wl_1_34
* pin wl_1_33
* pin wl_1_45
* pin wl_0_33
* pin wl_1_32
* pin wl_1_46
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_capped_replica_bitcell_array_0 1 2 3
+ 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31
+ 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57
+ 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106
+ 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125
+ 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144
+ 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239
+ 240 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258
+ 259 260
* net 1 wl_1_9
* net 2 wl_1_20
* net 3 wl_1_19
* net 4 wl_0_9
* net 5 wl_1_23
* net 6 wl_0_19
* net 7 wl_0_8
* net 8 wl_0_18
* net 9 wl_1_8
* net 10 wl_1_18
* net 11 wl_1_12
* net 12 wl_0_12
* net 13 wl_0_23
* net 14 wl_1_3
* net 15 wl_1_10
* net 16 wl_0_20
* net 17 wl_0_10
* net 18 wl_0_21
* net 19 wl_1_15
* net 20 wl_0_22
* net 21 wl_0_11
* net 22 wl_1_21
* net 23 wl_1_11
* net 24 wl_1_22
* net 25 wl_1_2
* net 26 wl_1_16
* net 27 wl_1_5
* net 28 wl_1_0
* net 29 wl_0_5
* net 30 wl_0_0
* net 31 wl_0_1
* net 32 wl_1_1
* net 33 wl_0_14
* net 34 wl_0_15
* net 35 wl_0_4
* net 36 wl_0_2
* net 37 wl_1_4
* net 38 wl_1_13
* net 39 wl_0_3
* net 40 wl_0_13
* net 41 wl_0_16
* net 42 wl_1_7
* net 43 wl_1_14
* net 44 wl_0_7
* net 45 wl_1_6
* net 46 rbl_wl_0_0
* net 47 wl_0_6
* net 48 wl_0_17
* net 49 wl_1_17
* net 50 bl_0_0
* net 51 bl_1_0
* net 52 br_1_0
* net 53 br_0_0
* net 54 bl_0_1
* net 55 bl_1_1
* net 56 br_1_1
* net 57 br_0_1
* net 58 bl_0_2
* net 59 bl_1_2
* net 60 br_1_2
* net 61 br_0_2
* net 62 bl_0_3
* net 63 bl_1_3
* net 64 br_1_3
* net 65 br_0_3
* net 66 bl_0_4
* net 67 bl_1_4
* net 68 br_1_4
* net 69 br_0_4
* net 70 bl_0_5
* net 71 bl_1_5
* net 72 br_1_5
* net 73 br_0_5
* net 74 bl_0_6
* net 75 bl_1_6
* net 76 br_1_6
* net 77 br_0_6
* net 78 bl_0_7
* net 79 bl_1_7
* net 80 br_1_7
* net 81 br_0_7
* net 82 bl_0_8
* net 83 bl_1_8
* net 84 br_1_8
* net 85 br_0_8
* net 86 bl_0_9
* net 87 bl_1_9
* net 88 br_1_9
* net 89 br_0_9
* net 90 bl_0_10
* net 91 bl_1_10
* net 92 br_1_10
* net 93 br_0_10
* net 94 bl_0_11
* net 95 bl_1_11
* net 96 br_1_11
* net 97 br_0_11
* net 98 bl_0_12
* net 99 bl_1_12
* net 100 br_1_12
* net 101 br_0_12
* net 102 bl_0_13
* net 103 bl_1_13
* net 104 br_1_13
* net 105 br_0_13
* net 106 bl_0_14
* net 107 bl_1_14
* net 108 br_1_14
* net 109 br_0_14
* net 110 bl_0_15
* net 111 bl_1_15
* net 112 br_1_15
* net 113 br_0_15
* net 114 wl_0_27
* net 115 wl_0_30
* net 116 wl_1_30
* net 117 wl_1_24
* net 118 wl_1_29
* net 119 wl_0_24
* net 120 wl_0_29
* net 121 wl_0_25
* net 122 wl_0_31
* net 123 wl_1_25
* net 124 wl_1_31
* net 125 wl_1_26
* net 126 wl_0_28
* net 127 wl_0_26
* net 128 wl_1_28
* net 129 wl_1_27
* net 130 bl_0_16
* net 131 bl_1_16
* net 132 br_1_16
* net 133 br_0_16
* net 134 bl_0_17
* net 135 bl_1_17
* net 136 br_1_17
* net 137 br_0_17
* net 138 bl_0_18
* net 139 bl_1_18
* net 140 br_1_18
* net 141 br_0_18
* net 142 bl_0_19
* net 143 bl_1_19
* net 144 br_1_19
* net 145 br_0_19
* net 146 bl_0_20
* net 147 bl_1_20
* net 148 br_1_20
* net 149 br_0_20
* net 150 bl_0_21
* net 151 bl_1_21
* net 152 br_1_21
* net 153 br_0_21
* net 154 bl_0_22
* net 155 bl_1_22
* net 156 br_1_22
* net 157 br_0_22
* net 158 bl_0_23
* net 159 bl_1_23
* net 160 br_1_23
* net 161 br_0_23
* net 162 bl_0_24
* net 163 bl_1_24
* net 164 br_1_24
* net 165 br_0_24
* net 166 bl_0_25
* net 167 bl_1_25
* net 168 br_1_25
* net 169 br_0_25
* net 170 bl_0_26
* net 171 bl_1_26
* net 172 br_1_26
* net 173 br_0_26
* net 174 bl_0_27
* net 175 bl_1_27
* net 176 br_1_27
* net 177 br_0_27
* net 178 bl_0_28
* net 179 bl_1_28
* net 180 br_1_28
* net 181 br_0_28
* net 182 bl_0_29
* net 183 bl_1_29
* net 184 br_1_29
* net 185 br_0_29
* net 186 bl_0_30
* net 187 bl_1_30
* net 188 br_1_30
* net 189 br_0_30
* net 190 bl_0_31
* net 191 bl_1_31
* net 192 br_1_31
* net 193 br_0_31
* net 194 wl_1_62
* net 195 wl_0_62
* net 196 rbl_wl_1_1
* net 197 wl_1_49
* net 198 wl_0_49
* net 199 wl_0_48
* net 200 wl_1_48
* net 201 wl_0_63
* net 202 wl_1_50
* net 203 wl_1_63
* net 204 wl_1_47
* net 205 wl_0_50
* net 206 wl_0_47
* net 207 wl_0_59
* net 208 wl_1_55
* net 209 wl_0_58
* net 210 wl_1_58
* net 211 wl_1_59
* net 212 wl_0_32
* net 213 wl_1_57
* net 214 wl_0_57
* net 215 wl_1_60
* net 216 wl_0_56
* net 217 wl_1_56
* net 218 wl_0_60
* net 219 wl_0_51
* net 220 wl_0_55
* net 221 wl_0_61
* net 222 wl_0_54
* net 223 wl_1_54
* net 224 wl_1_53
* net 225 wl_0_53
* net 226 wl_0_52
* net 227 wl_1_52
* net 228 wl_1_51
* net 229 wl_1_61
* net 230 wl_0_39
* net 231 wl_0_44
* net 232 wl_0_35
* net 233 wl_1_35
* net 234 wl_1_36
* net 235 wl_1_44
* net 236 wl_0_36
* net 237 wl_0_37
* net 238 wl_1_37
* net 239 wl_1_38
* net 240 wl_0_38
* net 241 wl_0_46
* net 242 wl_1_39
* net 243 wl_1_43
* net 244 wl_1_40
* net 245 wl_0_40
* net 246 wl_0_43
* net 247 wl_0_41
* net 248 wl_1_41
* net 249 wl_1_42
* net 250 wl_0_42
* net 251 wl_0_45
* net 252 wl_0_34
* net 253 wl_1_34
* net 254 wl_1_33
* net 255 wl_1_45
* net 256 wl_0_33
* net 257 wl_1_32
* net 258 wl_1_46
* net 259 vdd
* net 260 gnd
* cell instance $1 r0 *1 0.935,0.25
X$1 260 260 46 260 28 30 31 32 25 36 39 14 37 35 29 27 45 47 44 42 9 7 4 1 15
+ 17 21 23 11 12 40 38 43 33 34 19 26 41 48 49 10 8 6 3 2 16 18 22 24 20 13 5
+ 117 119 121 123 125 127 114 129 128 126 120 118 116 115 122 124 257 212 256
+ 254 253 252 232 233 234 236 237 238 239 240 230 242 244 245 247 248 249 250
+ 246 243 235 231 251 255 258 241 206 204 200 199 198 197 202 205 219 228 227
+ 226 225 224 223 222 220 208 217 216 214 213 210 209 207 211 215 218 221 229
+ 194 195 201 203 196 260 260 260 259 260
+ custom_sram_1r1w_32_256_freepdk45_dummy_array_2
* cell instance $2 r0 *1 2.11,1.745
X$2 46 260 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72
+ 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98
+ 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 130 131 132 133
+ 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152
+ 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171
+ 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190
+ 191 192 193 28 30 31 32 36 25 14 39 35 37 27 29 45 47 42 44 9 7 1 4 15 17 21
+ 23 12 11 38 40 33 43 34 19 41 26 49 48 10 8 3 6 2 16 18 22 24 20 13 5 117 119
+ 123 121 127 125 129 114 128 126 118 120 116 115 124 122 257 212 256 254 252
+ 253 233 232 236 234 238 237 240 239 242 230 245 244 248 247 250 249 243 246
+ 235 231 255 251 258 241 204 206 200 199 197 198 205 202 228 219 226 227 225
+ 224 223 222 220 208 216 217 213 214 210 209 211 207 218 215 221 229 194 195
+ 203 201 260 196 259 260
+ custom_sram_1r1w_32_256_freepdk45_replica_bitcell_array_0
* cell instance $3 r0 *1 39.71,0.25
X$3 260 260 46 260 28 30 31 32 25 36 39 14 37 35 29 27 45 47 44 42 9 7 4 1 15
+ 17 21 23 11 12 40 38 43 33 34 19 26 41 48 49 10 8 6 3 2 16 18 22 24 20 13 5
+ 117 119 121 123 125 127 114 129 128 126 120 118 116 115 122 124 257 212 256
+ 254 253 252 232 233 234 236 237 238 239 240 230 242 244 245 247 248 249 250
+ 246 243 235 231 251 255 258 241 206 204 200 199 198 197 202 205 219 228 227
+ 226 225 224 223 222 220 208 217 216 214 213 210 209 207 211 215 218 221 229
+ 194 195 201 203 196 260 260 260 259 260
+ custom_sram_1r1w_32_256_freepdk45_dummy_array_7
* cell instance $4 r0 *1 2.11,0.25
X$4 260 260 259 260 custom_sram_1r1w_32_256_freepdk45_dummy_array_6
* cell instance $5 m0 *1 2.11,101.91
X$5 260 260 259 260 custom_sram_1r1w_32_256_freepdk45_dummy_array_5
.ENDS custom_sram_1r1w_32_256_freepdk45_capped_replica_bitcell_array_0

* cell custom_sram_1r1w_32_256_freepdk45_capped_replica_bitcell_array
* pin wl_1_9
* pin wl_0_23
* pin rbl_wl_0_0
* pin wl_0_16
* pin wl_0_17
* pin wl_1_19
* pin wl_1_23
* pin wl_0_9
* pin wl_0_18
* pin wl_1_24
* pin wl_1_17
* pin wl_0_24
* pin wl_0_19
* pin wl_0_20
* pin wl_1_11
* pin wl_1_14
* pin wl_0_14
* pin wl_1_13
* pin wl_0_13
* pin wl_0_12
* pin wl_1_12
* pin wl_1_18
* pin wl_0_15
* pin wl_1_15
* pin wl_0_22
* pin wl_0_11
* pin wl_0_10
* pin wl_0_21
* pin wl_1_10
* pin wl_1_21
* pin wl_1_20
* pin wl_1_16
* pin wl_1_22
* pin wl_0_8
* pin wl_1_0
* pin wl_0_0
* pin wl_0_1
* pin wl_1_1
* pin wl_1_2
* pin wl_0_2
* pin wl_0_3
* pin wl_1_3
* pin wl_1_4
* pin wl_0_4
* pin wl_0_5
* pin wl_1_8
* pin wl_1_7
* pin wl_0_7
* pin wl_0_6
* pin wl_1_6
* pin wl_1_5
* pin rbl_bl_0_0
* pin rbl_bl_1_0
* pin rbl_br_1_0
* pin rbl_br_0_0
* pin bl_0_0
* pin bl_1_0
* pin br_1_0
* pin br_0_0
* pin bl_0_1
* pin bl_1_1
* pin br_1_1
* pin br_0_1
* pin bl_0_2
* pin bl_1_2
* pin br_1_2
* pin br_0_2
* pin bl_0_3
* pin bl_1_3
* pin br_1_3
* pin br_0_3
* pin bl_0_4
* pin bl_1_4
* pin br_1_4
* pin br_0_4
* pin bl_0_5
* pin bl_1_5
* pin br_1_5
* pin br_0_5
* pin bl_0_6
* pin bl_1_6
* pin br_1_6
* pin br_0_6
* pin bl_0_7
* pin bl_1_7
* pin br_1_7
* pin br_0_7
* pin bl_0_8
* pin bl_1_8
* pin br_1_8
* pin br_0_8
* pin bl_0_9
* pin bl_1_9
* pin br_1_9
* pin br_0_9
* pin bl_0_10
* pin bl_1_10
* pin br_1_10
* pin br_0_10
* pin bl_0_11
* pin bl_1_11
* pin br_1_11
* pin br_0_11
* pin bl_0_12
* pin bl_1_12
* pin br_1_12
* pin br_0_12
* pin bl_0_13
* pin bl_1_13
* pin br_1_13
* pin br_0_13
* pin bl_0_14
* pin bl_1_14
* pin br_1_14
* pin br_0_14
* pin bl_0_15
* pin bl_1_15
* pin wl_1_31
* pin wl_1_30
* pin wl_0_30
* pin wl_0_31
* pin wl_0_29
* pin wl_0_28
* pin wl_1_28
* pin wl_1_27
* pin wl_0_27
* pin wl_0_25
* pin wl_0_26
* pin wl_1_29
* pin wl_1_26
* pin wl_1_25
* pin br_1_15
* pin br_0_15
* pin bl_0_16
* pin bl_1_16
* pin br_1_16
* pin br_0_16
* pin bl_0_17
* pin bl_1_17
* pin br_1_17
* pin br_0_17
* pin bl_0_18
* pin bl_1_18
* pin br_1_18
* pin br_0_18
* pin bl_0_19
* pin bl_1_19
* pin br_1_19
* pin br_0_19
* pin bl_0_20
* pin bl_1_20
* pin br_1_20
* pin br_0_20
* pin bl_0_21
* pin bl_1_21
* pin br_1_21
* pin br_0_21
* pin bl_0_22
* pin bl_1_22
* pin br_1_22
* pin br_0_22
* pin bl_0_23
* pin bl_1_23
* pin br_1_23
* pin br_0_23
* pin bl_0_24
* pin bl_1_24
* pin br_1_24
* pin br_0_24
* pin bl_0_25
* pin bl_1_25
* pin br_1_25
* pin br_0_25
* pin bl_0_26
* pin bl_1_26
* pin br_1_26
* pin br_0_26
* pin bl_0_27
* pin bl_1_27
* pin br_1_27
* pin br_0_27
* pin bl_0_28
* pin bl_1_28
* pin br_1_28
* pin br_0_28
* pin bl_0_29
* pin bl_1_29
* pin br_1_29
* pin br_0_29
* pin bl_0_30
* pin bl_1_30
* pin br_1_30
* pin br_0_30
* pin bl_0_31
* pin bl_1_31
* pin br_1_31
* pin br_0_31
* pin wl_0_47
* pin wl_1_52
* pin rbl_wl_1_1
* pin wl_1_51
* pin wl_1_56
* pin wl_1_48
* pin wl_0_46
* pin wl_0_56
* pin wl_1_46
* pin wl_0_52
* pin wl_0_45
* pin wl_0_49
* pin wl_0_53
* pin wl_0_33
* pin wl_1_53
* pin wl_0_50
* pin wl_1_50
* pin wl_1_54
* pin wl_0_51
* pin wl_1_49
* pin wl_1_47
* pin wl_0_54
* pin wl_0_60
* pin wl_1_34
* pin wl_0_48
* pin wl_0_55
* pin wl_1_55
* pin wl_0_34
* pin wl_1_60
* pin wl_1_57
* pin wl_1_59
* pin wl_1_42
* pin wl_0_59
* pin wl_1_36
* pin wl_0_62
* pin wl_0_36
* pin wl_1_41
* pin wl_1_45
* pin wl_0_41
* pin wl_0_32
* pin wl_1_62
* pin wl_0_40
* pin wl_1_40
* pin wl_0_58
* pin wl_1_39
* pin wl_0_39
* pin wl_0_37
* pin wl_1_37
* pin wl_0_38
* pin wl_1_38
* pin wl_1_32
* pin wl_0_61
* pin wl_1_58
* pin wl_0_42
* pin wl_0_44
* pin wl_1_44
* pin wl_0_35
* pin wl_1_43
* pin wl_1_63
* pin wl_0_43
* pin wl_1_33
* pin wl_1_61
* pin wl_0_57
* pin wl_0_63
* pin wl_1_35
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_capped_replica_bitcell_array 1 2 3 4
+ 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31
+ 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57
+ 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106
+ 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125
+ 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144
+ 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239
+ 240 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258
+ 259 260 261 262 263 264
* net 1 wl_1_9
* net 2 wl_0_23
* net 3 rbl_wl_0_0
* net 4 wl_0_16
* net 5 wl_0_17
* net 6 wl_1_19
* net 7 wl_1_23
* net 8 wl_0_9
* net 9 wl_0_18
* net 10 wl_1_24
* net 11 wl_1_17
* net 12 wl_0_24
* net 13 wl_0_19
* net 14 wl_0_20
* net 15 wl_1_11
* net 16 wl_1_14
* net 17 wl_0_14
* net 18 wl_1_13
* net 19 wl_0_13
* net 20 wl_0_12
* net 21 wl_1_12
* net 22 wl_1_18
* net 23 wl_0_15
* net 24 wl_1_15
* net 25 wl_0_22
* net 26 wl_0_11
* net 27 wl_0_10
* net 28 wl_0_21
* net 29 wl_1_10
* net 30 wl_1_21
* net 31 wl_1_20
* net 32 wl_1_16
* net 33 wl_1_22
* net 34 wl_0_8
* net 35 wl_1_0
* net 36 wl_0_0
* net 37 wl_0_1
* net 38 wl_1_1
* net 39 wl_1_2
* net 40 wl_0_2
* net 41 wl_0_3
* net 42 wl_1_3
* net 43 wl_1_4
* net 44 wl_0_4
* net 45 wl_0_5
* net 46 wl_1_8
* net 47 wl_1_7
* net 48 wl_0_7
* net 49 wl_0_6
* net 50 wl_1_6
* net 51 wl_1_5
* net 52 rbl_bl_0_0
* net 53 rbl_bl_1_0
* net 54 rbl_br_1_0
* net 55 rbl_br_0_0
* net 56 bl_0_0
* net 57 bl_1_0
* net 58 br_1_0
* net 59 br_0_0
* net 60 bl_0_1
* net 61 bl_1_1
* net 62 br_1_1
* net 63 br_0_1
* net 64 bl_0_2
* net 65 bl_1_2
* net 66 br_1_2
* net 67 br_0_2
* net 68 bl_0_3
* net 69 bl_1_3
* net 70 br_1_3
* net 71 br_0_3
* net 72 bl_0_4
* net 73 bl_1_4
* net 74 br_1_4
* net 75 br_0_4
* net 76 bl_0_5
* net 77 bl_1_5
* net 78 br_1_5
* net 79 br_0_5
* net 80 bl_0_6
* net 81 bl_1_6
* net 82 br_1_6
* net 83 br_0_6
* net 84 bl_0_7
* net 85 bl_1_7
* net 86 br_1_7
* net 87 br_0_7
* net 88 bl_0_8
* net 89 bl_1_8
* net 90 br_1_8
* net 91 br_0_8
* net 92 bl_0_9
* net 93 bl_1_9
* net 94 br_1_9
* net 95 br_0_9
* net 96 bl_0_10
* net 97 bl_1_10
* net 98 br_1_10
* net 99 br_0_10
* net 100 bl_0_11
* net 101 bl_1_11
* net 102 br_1_11
* net 103 br_0_11
* net 104 bl_0_12
* net 105 bl_1_12
* net 106 br_1_12
* net 107 br_0_12
* net 108 bl_0_13
* net 109 bl_1_13
* net 110 br_1_13
* net 111 br_0_13
* net 112 bl_0_14
* net 113 bl_1_14
* net 114 br_1_14
* net 115 br_0_14
* net 116 bl_0_15
* net 117 bl_1_15
* net 118 wl_1_31
* net 119 wl_1_30
* net 120 wl_0_30
* net 121 wl_0_31
* net 122 wl_0_29
* net 123 wl_0_28
* net 124 wl_1_28
* net 125 wl_1_27
* net 126 wl_0_27
* net 127 wl_0_25
* net 128 wl_0_26
* net 129 wl_1_29
* net 130 wl_1_26
* net 131 wl_1_25
* net 132 br_1_15
* net 133 br_0_15
* net 134 bl_0_16
* net 135 bl_1_16
* net 136 br_1_16
* net 137 br_0_16
* net 138 bl_0_17
* net 139 bl_1_17
* net 140 br_1_17
* net 141 br_0_17
* net 142 bl_0_18
* net 143 bl_1_18
* net 144 br_1_18
* net 145 br_0_18
* net 146 bl_0_19
* net 147 bl_1_19
* net 148 br_1_19
* net 149 br_0_19
* net 150 bl_0_20
* net 151 bl_1_20
* net 152 br_1_20
* net 153 br_0_20
* net 154 bl_0_21
* net 155 bl_1_21
* net 156 br_1_21
* net 157 br_0_21
* net 158 bl_0_22
* net 159 bl_1_22
* net 160 br_1_22
* net 161 br_0_22
* net 162 bl_0_23
* net 163 bl_1_23
* net 164 br_1_23
* net 165 br_0_23
* net 166 bl_0_24
* net 167 bl_1_24
* net 168 br_1_24
* net 169 br_0_24
* net 170 bl_0_25
* net 171 bl_1_25
* net 172 br_1_25
* net 173 br_0_25
* net 174 bl_0_26
* net 175 bl_1_26
* net 176 br_1_26
* net 177 br_0_26
* net 178 bl_0_27
* net 179 bl_1_27
* net 180 br_1_27
* net 181 br_0_27
* net 182 bl_0_28
* net 183 bl_1_28
* net 184 br_1_28
* net 185 br_0_28
* net 186 bl_0_29
* net 187 bl_1_29
* net 188 br_1_29
* net 189 br_0_29
* net 190 bl_0_30
* net 191 bl_1_30
* net 192 br_1_30
* net 193 br_0_30
* net 194 bl_0_31
* net 195 bl_1_31
* net 196 br_1_31
* net 197 br_0_31
* net 198 wl_0_47
* net 199 wl_1_52
* net 200 rbl_wl_1_1
* net 201 wl_1_51
* net 202 wl_1_56
* net 203 wl_1_48
* net 204 wl_0_46
* net 205 wl_0_56
* net 206 wl_1_46
* net 207 wl_0_52
* net 208 wl_0_45
* net 209 wl_0_49
* net 210 wl_0_53
* net 211 wl_0_33
* net 212 wl_1_53
* net 213 wl_0_50
* net 214 wl_1_50
* net 215 wl_1_54
* net 216 wl_0_51
* net 217 wl_1_49
* net 218 wl_1_47
* net 219 wl_0_54
* net 220 wl_0_60
* net 221 wl_1_34
* net 222 wl_0_48
* net 223 wl_0_55
* net 224 wl_1_55
* net 225 wl_0_34
* net 226 wl_1_60
* net 227 wl_1_57
* net 228 wl_1_59
* net 229 wl_1_42
* net 230 wl_0_59
* net 231 wl_1_36
* net 232 wl_0_62
* net 233 wl_0_36
* net 234 wl_1_41
* net 235 wl_1_45
* net 236 wl_0_41
* net 237 wl_0_32
* net 238 wl_1_62
* net 239 wl_0_40
* net 240 wl_1_40
* net 241 wl_0_58
* net 242 wl_1_39
* net 243 wl_0_39
* net 244 wl_0_37
* net 245 wl_1_37
* net 246 wl_0_38
* net 247 wl_1_38
* net 248 wl_1_32
* net 249 wl_0_61
* net 250 wl_1_58
* net 251 wl_0_42
* net 252 wl_0_44
* net 253 wl_1_44
* net 254 wl_0_35
* net 255 wl_1_43
* net 256 wl_1_63
* net 257 wl_0_43
* net 258 wl_1_33
* net 259 wl_1_61
* net 260 wl_0_57
* net 261 wl_0_63
* net 262 wl_1_35
* net 263 vdd
* net 264 gnd
* cell instance $1 r0 *1 0.935,0.25
X$1 264 264 3 264 35 36 37 38 39 40 41 42 43 44 45 51 50 49 48 47 46 34 8 1 29
+ 27 26 15 21 20 19 18 16 17 23 24 32 4 5 11 22 9 13 6 31 14 28 30 33 25 2 7 10
+ 12 127 131 130 128 126 125 124 123 122 129 119 120 121 118 248 237 211 258
+ 221 225 254 262 231 233 244 245 247 246 243 242 240 239 236 234 229 251 257
+ 255 253 252 208 235 206 204 198 218 203 222 209 217 214 213 216 201 199 207
+ 210 212 215 219 223 224 202 205 260 227 250 241 230 228 226 220 249 259 238
+ 232 261 256 200 264 264 264 263 264
+ custom_sram_1r1w_32_256_freepdk45_dummy_array_2
* cell instance $2 r0 *1 2.11,1.745
X$2 3 264 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74
+ 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99
+ 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 132
+ 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151
+ 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170
+ 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189
+ 190 191 192 193 194 195 196 197 35 36 38 37 40 39 42 41 44 43 51 45 49 50 48
+ 47 34 46 8 1 27 29 15 26 20 21 18 19 17 16 24 23 4 32 11 5 9 22 6 13 14 31 30
+ 28 33 25 2 7 10 12 131 127 128 130 125 126 123 124 129 122 120 119 118 121
+ 248 237 258 211 225 221 262 254 233 231 244 245 246 247 243 242 239 240 234
+ 236 251 229 255 257 252 253 235 208 204 206 218 198 222 203 209 217 213 214
+ 201 216 207 199 212 210 215 219 224 223 202 205 227 260 250 241 228 230 220
+ 226 249 259 238 232 261 256 200 264 263 264
+ custom_sram_1r1w_32_256_freepdk45_replica_bitcell_array
* cell instance $3 r0 *1 40.885,0.25
X$3 264 264 3 264 35 36 37 38 39 40 41 42 43 44 45 51 50 49 48 47 46 34 8 1 29
+ 27 26 15 21 20 19 18 16 17 23 24 32 4 5 11 22 9 13 6 31 14 28 30 33 25 2 7 10
+ 12 127 131 130 128 126 125 124 123 122 129 119 120 121 118 248 237 211 258
+ 221 225 254 262 231 233 244 245 247 246 243 242 240 239 236 234 229 251 257
+ 255 253 252 208 235 206 204 198 218 203 222 209 217 214 213 216 201 199 207
+ 210 212 215 219 223 224 202 205 260 227 250 241 230 228 226 220 249 259 238
+ 232 261 256 200 264 264 264 263 264
+ custom_sram_1r1w_32_256_freepdk45_dummy_array_3
* cell instance $4 r0 *1 2.11,0.25
X$4 264 264 263 264 custom_sram_1r1w_32_256_freepdk45_dummy_array_1
* cell instance $5 m0 *1 2.11,101.91
X$5 264 264 263 264 custom_sram_1r1w_32_256_freepdk45_dummy_array_0
.ENDS custom_sram_1r1w_32_256_freepdk45_capped_replica_bitcell_array

* cell custom_sram_1r1w_32_256_freepdk45_wordline_buffer_array
* pin in_0
* pin out_0
* pin in_1
* pin out_1
* pin in_2
* pin out_2
* pin in_3
* pin out_3
* pin in_4
* pin out_4
* pin in_5
* pin out_5
* pin in_6
* pin out_6
* pin in_7
* pin out_7
* pin in_8
* pin out_8
* pin in_9
* pin out_9
* pin in_10
* pin out_10
* pin in_11
* pin out_11
* pin in_12
* pin out_12
* pin in_13
* pin out_13
* pin in_14
* pin out_14
* pin in_15
* pin out_15
* pin in_16
* pin out_16
* pin in_17
* pin out_17
* pin in_18
* pin out_18
* pin in_19
* pin out_19
* pin in_20
* pin out_20
* pin in_21
* pin out_21
* pin in_22
* pin out_22
* pin in_23
* pin out_23
* pin in_24
* pin out_24
* pin in_25
* pin out_25
* pin in_26
* pin out_26
* pin in_27
* pin out_27
* pin in_28
* pin out_28
* pin in_29
* pin out_29
* pin in_30
* pin out_30
* pin in_31
* pin out_31
* pin in_32
* pin out_32
* pin in_33
* pin out_33
* pin in_34
* pin out_34
* pin in_35
* pin out_35
* pin in_36
* pin out_36
* pin in_37
* pin out_37
* pin in_38
* pin out_38
* pin in_39
* pin out_39
* pin in_40
* pin out_40
* pin in_41
* pin out_41
* pin in_42
* pin out_42
* pin in_43
* pin out_43
* pin in_44
* pin out_44
* pin in_45
* pin out_45
* pin in_46
* pin out_46
* pin in_47
* pin out_47
* pin in_48
* pin out_48
* pin in_49
* pin out_49
* pin in_50
* pin out_50
* pin in_51
* pin out_51
* pin in_52
* pin out_52
* pin in_53
* pin out_53
* pin in_54
* pin out_54
* pin in_55
* pin out_55
* pin in_56
* pin out_56
* pin in_57
* pin out_57
* pin in_58
* pin out_58
* pin in_59
* pin out_59
* pin in_60
* pin out_60
* pin in_61
* pin out_61
* pin in_62
* pin out_62
* pin in_63
* pin out_63
* pin in_64
* pin out_64
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_wordline_buffer_array 1 2 3 4 5 6 7 8
+ 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34
+ 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86
+ 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108
+ 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127
+ 128 129 130 131 132
* net 1 in_0
* net 2 out_0
* net 3 in_1
* net 4 out_1
* net 5 in_2
* net 6 out_2
* net 7 in_3
* net 8 out_3
* net 9 in_4
* net 10 out_4
* net 11 in_5
* net 12 out_5
* net 13 in_6
* net 14 out_6
* net 15 in_7
* net 16 out_7
* net 17 in_8
* net 18 out_8
* net 19 in_9
* net 20 out_9
* net 21 in_10
* net 22 out_10
* net 23 in_11
* net 24 out_11
* net 25 in_12
* net 26 out_12
* net 27 in_13
* net 28 out_13
* net 29 in_14
* net 30 out_14
* net 31 in_15
* net 32 out_15
* net 33 in_16
* net 34 out_16
* net 35 in_17
* net 36 out_17
* net 37 in_18
* net 38 out_18
* net 39 in_19
* net 40 out_19
* net 41 in_20
* net 42 out_20
* net 43 in_21
* net 44 out_21
* net 45 in_22
* net 46 out_22
* net 47 in_23
* net 48 out_23
* net 49 in_24
* net 50 out_24
* net 51 in_25
* net 52 out_25
* net 53 in_26
* net 54 out_26
* net 55 in_27
* net 56 out_27
* net 57 in_28
* net 58 out_28
* net 59 in_29
* net 60 out_29
* net 61 in_30
* net 62 out_30
* net 63 in_31
* net 64 out_31
* net 65 in_32
* net 66 out_32
* net 67 in_33
* net 68 out_33
* net 69 in_34
* net 70 out_34
* net 71 in_35
* net 72 out_35
* net 73 in_36
* net 74 out_36
* net 75 in_37
* net 76 out_37
* net 77 in_38
* net 78 out_38
* net 79 in_39
* net 80 out_39
* net 81 in_40
* net 82 out_40
* net 83 in_41
* net 84 out_41
* net 85 in_42
* net 86 out_42
* net 87 in_43
* net 88 out_43
* net 89 in_44
* net 90 out_44
* net 91 in_45
* net 92 out_45
* net 93 in_46
* net 94 out_46
* net 95 in_47
* net 96 out_47
* net 97 in_48
* net 98 out_48
* net 99 in_49
* net 100 out_49
* net 101 in_50
* net 102 out_50
* net 103 in_51
* net 104 out_51
* net 105 in_52
* net 106 out_52
* net 107 in_53
* net 108 out_53
* net 109 in_54
* net 110 out_54
* net 111 in_55
* net 112 out_55
* net 113 in_56
* net 114 out_56
* net 115 in_57
* net 116 out_57
* net 117 in_58
* net 118 out_58
* net 119 in_59
* net 120 out_59
* net 121 in_60
* net 122 out_60
* net 123 in_61
* net 124 out_61
* net 125 in_62
* net 126 out_62
* net 127 in_63
* net 128 out_63
* net 129 in_64
* net 130 out_64
* net 131 vdd
* net 132 gnd
* cell instance $1 m0 *1 0,1.495
X$1 1 2 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $2 r0 *1 0,1.495
X$2 3 4 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $3 m0 *1 0,4.485
X$3 5 6 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $4 r0 *1 0,4.485
X$4 7 8 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $5 m0 *1 0,7.475
X$5 9 10 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $6 r0 *1 0,7.475
X$6 11 12 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $7 m0 *1 0,10.465
X$7 13 14 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $8 r0 *1 0,10.465
X$8 15 16 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $9 m0 *1 0,13.455
X$9 17 18 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $10 r0 *1 0,13.455
X$10 19 20 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $11 m0 *1 0,16.445
X$11 21 22 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $12 r0 *1 0,16.445
X$12 23 24 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $13 m0 *1 0,19.435
X$13 25 26 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $14 r0 *1 0,19.435
X$14 27 28 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $15 m0 *1 0,22.425
X$15 29 30 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $16 r0 *1 0,22.425
X$16 31 32 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $17 m0 *1 0,25.415
X$17 33 34 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $18 r0 *1 0,25.415
X$18 35 36 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $19 m0 *1 0,28.405
X$19 37 38 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $20 r0 *1 0,28.405
X$20 39 40 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $21 m0 *1 0,31.395
X$21 41 42 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $22 r0 *1 0,31.395
X$22 43 44 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $23 m0 *1 0,34.385
X$23 45 46 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $24 r0 *1 0,34.385
X$24 47 48 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $25 m0 *1 0,37.375
X$25 49 50 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $26 r0 *1 0,37.375
X$26 51 52 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $27 m0 *1 0,40.365
X$27 53 54 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $28 r0 *1 0,40.365
X$28 55 56 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $29 m0 *1 0,43.355
X$29 57 58 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $30 r0 *1 0,43.355
X$30 59 60 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $31 m0 *1 0,46.345
X$31 61 62 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $32 r0 *1 0,46.345
X$32 63 64 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $33 m0 *1 0,49.335
X$33 65 66 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $34 r0 *1 0,49.335
X$34 67 68 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $35 m0 *1 0,52.325
X$35 69 70 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $36 r0 *1 0,52.325
X$36 71 72 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $37 m0 *1 0,55.315
X$37 73 74 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $38 r0 *1 0,55.315
X$38 75 76 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $39 m0 *1 0,58.305
X$39 77 78 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $40 r0 *1 0,58.305
X$40 79 80 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $41 m0 *1 0,61.295
X$41 81 82 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $42 r0 *1 0,61.295
X$42 83 84 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $43 m0 *1 0,64.285
X$43 85 86 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $44 r0 *1 0,64.285
X$44 87 88 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $45 m0 *1 0,67.275
X$45 89 90 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $46 r0 *1 0,67.275
X$46 91 92 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $47 m0 *1 0,70.265
X$47 93 94 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $48 r0 *1 0,70.265
X$48 95 96 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $49 m0 *1 0,73.255
X$49 97 98 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $50 r0 *1 0,73.255
X$50 99 100 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $51 m0 *1 0,76.245
X$51 101 102 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $52 r0 *1 0,76.245
X$52 103 104 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $53 m0 *1 0,79.235
X$53 105 106 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $54 r0 *1 0,79.235
X$54 107 108 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $55 m0 *1 0,82.225
X$55 109 110 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $56 r0 *1 0,82.225
X$56 111 112 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $57 m0 *1 0,85.215
X$57 113 114 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $58 r0 *1 0,85.215
X$58 115 116 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $59 m0 *1 0,88.205
X$59 117 118 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $60 r0 *1 0,88.205
X$60 119 120 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $61 m0 *1 0,91.195
X$61 121 122 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $62 r0 *1 0,91.195
X$62 123 124 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $63 m0 *1 0,94.185
X$63 125 126 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $64 r0 *1 0,94.185
X$64 127 128 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
* cell instance $65 m0 *1 0,97.175
X$65 129 130 131 132 custom_sram_1r1w_32_256_freepdk45_pinv
.ENDS custom_sram_1r1w_32_256_freepdk45_wordline_buffer_array

* cell custom_sram_1r1w_32_256_freepdk45_pdriver
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pdriver 1 2 3 4
* net 1 Z
* net 2 A
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 custom_sram_1r1w_32_256_freepdk45_pinv_3
.ENDS custom_sram_1r1w_32_256_freepdk45_pdriver

* cell custom_sram_1r1w_32_256_freepdk45_pnand2_0
* pin A
* pin B
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pnand2_0 1 2 3 4 5
* net 1 A
* net 2 B
* net 3 Z
* net 4 vdd
* net 5 gnd
* device instance $1 r0 *1 0.2325,2.21 PMOS_VTG
M$1 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,2.21 PMOS_VTG
M$2 3 2 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.2325,0.215 NMOS_VTG
M$3 5 1 6 5 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $4 r0 *1 0.4475,0.215 NMOS_VTG
M$4 6 2 3 5 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS custom_sram_1r1w_32_256_freepdk45_pnand2_0

* cell custom_sram_1r1w_32_256_freepdk45_pbuf
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pbuf 2 3 4 5
* net 2 Z
* net 3 A
* net 4 vdd
* net 5 gnd
* cell instance $1 r0 *1 0,0
X$1 3 1 4 5 custom_sram_1r1w_32_256_freepdk45_pinv_0
* cell instance $2 r0 *1 0.6875,0
X$2 1 2 4 5 custom_sram_1r1w_32_256_freepdk45_pinv_1
.ENDS custom_sram_1r1w_32_256_freepdk45_pbuf

* cell custom_sram_1r1w_32_256_freepdk45_and2_dec
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_and2_dec 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0,0
X$1 3 4 1 5 6 custom_sram_1r1w_32_256_freepdk45_pnand2
* cell instance $2 r0 *1 0.9025,0
X$2 1 2 5 6 custom_sram_1r1w_32_256_freepdk45_pinv_0
.ENDS custom_sram_1r1w_32_256_freepdk45_and2_dec

* cell custom_sram_1r1w_32_256_freepdk45_pnand3
* pin A
* pin B
* pin C
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pnand3 1 2 3 4 5 6
* net 1 A
* net 2 B
* net 3 C
* net 4 Z
* net 5 vdd
* net 6 gnd
* device instance $1 r0 *1 0.2325,1.235 PMOS_VTG
M$1 5 1 4 5 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,1.235 PMOS_VTG
M$2 4 2 5 5 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.022275P PS=0.435U
+ PD=0.435U
* device instance $3 r0 *1 0.6625,1.235 PMOS_VTG
M$3 5 3 4 5 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $4 r0 *1 0.2325,0.215 NMOS_VTG
M$4 6 1 8 6 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $5 r0 *1 0.4475,0.215 NMOS_VTG
M$5 8 2 7 6 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.01485P PS=0.345U PD=0.345U
* device instance $6 r0 *1 0.6625,0.215 NMOS_VTG
M$6 7 3 4 6 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS custom_sram_1r1w_32_256_freepdk45_pnand3

* cell custom_sram_1r1w_32_256_freepdk45_replica_bitcell_array_1
* pin rbl_wl_0_1
* pin rbl_wl_0_0
* pin bl_0_0
* pin bl_1_0
* pin br_1_0
* pin br_0_0
* pin bl_0_1
* pin bl_1_1
* pin br_1_1
* pin br_0_1
* pin bl_0_2
* pin bl_1_2
* pin br_1_2
* pin br_0_2
* pin bl_0_3
* pin bl_1_3
* pin br_1_3
* pin br_0_3
* pin bl_0_4
* pin bl_1_4
* pin br_1_4
* pin br_0_4
* pin bl_0_5
* pin bl_1_5
* pin br_1_5
* pin br_0_5
* pin bl_0_6
* pin bl_1_6
* pin br_1_6
* pin br_0_6
* pin bl_0_7
* pin bl_1_7
* pin br_1_7
* pin br_0_7
* pin bl_0_8
* pin bl_1_8
* pin br_1_8
* pin br_0_8
* pin bl_0_9
* pin bl_1_9
* pin br_1_9
* pin br_0_9
* pin bl_0_10
* pin bl_1_10
* pin br_1_10
* pin br_0_10
* pin bl_0_11
* pin bl_1_11
* pin br_1_11
* pin br_0_11
* pin bl_0_12
* pin bl_1_12
* pin br_1_12
* pin br_0_12
* pin bl_0_13
* pin bl_1_13
* pin br_1_13
* pin br_0_13
* pin bl_0_14
* pin bl_1_14
* pin br_1_14
* pin br_0_14
* pin bl_0_15
* pin bl_1_15
* pin br_1_15
* pin br_0_15
* pin bl_0_16
* pin bl_1_16
* pin br_1_16
* pin br_0_16
* pin bl_0_17
* pin bl_1_17
* pin br_1_17
* pin br_0_17
* pin bl_0_18
* pin bl_1_18
* pin br_1_18
* pin br_0_18
* pin bl_0_19
* pin bl_1_19
* pin br_1_19
* pin br_0_19
* pin bl_0_20
* pin bl_1_20
* pin br_1_20
* pin br_0_20
* pin bl_0_21
* pin bl_1_21
* pin br_1_21
* pin br_0_21
* pin bl_0_22
* pin bl_1_22
* pin br_1_22
* pin br_0_22
* pin bl_0_23
* pin bl_1_23
* pin br_1_23
* pin br_0_23
* pin bl_0_24
* pin bl_1_24
* pin br_1_24
* pin br_0_24
* pin bl_0_25
* pin bl_1_25
* pin br_1_25
* pin br_0_25
* pin bl_0_26
* pin bl_1_26
* pin br_1_26
* pin br_0_26
* pin bl_0_27
* pin bl_1_27
* pin br_1_27
* pin br_0_27
* pin bl_0_28
* pin bl_1_28
* pin br_1_28
* pin br_0_28
* pin bl_0_29
* pin bl_1_29
* pin br_1_29
* pin br_0_29
* pin bl_0_30
* pin bl_1_30
* pin br_1_30
* pin br_0_30
* pin bl_0_31
* pin bl_1_31
* pin br_1_31
* pin br_0_31
* pin rbl_bl_0_1
* pin rbl_bl_1_1
* pin rbl_br_1_1
* pin rbl_br_0_1
* pin wl_0_0
* pin wl_1_0
* pin wl_1_1
* pin wl_0_1
* pin wl_1_2
* pin wl_0_2
* pin wl_1_3
* pin wl_0_3
* pin wl_1_4
* pin wl_0_4
* pin wl_1_5
* pin wl_0_5
* pin wl_0_6
* pin wl_1_6
* pin wl_1_7
* pin wl_0_7
* pin wl_0_8
* pin wl_1_8
* pin wl_1_9
* pin wl_0_9
* pin wl_1_10
* pin wl_0_10
* pin wl_1_11
* pin wl_0_11
* pin wl_1_12
* pin wl_0_12
* pin wl_1_13
* pin wl_0_13
* pin wl_0_14
* pin wl_1_14
* pin wl_1_15
* pin wl_0_15
* pin wl_0_16
* pin wl_1_16
* pin wl_1_17
* pin wl_0_17
* pin wl_0_18
* pin wl_1_18
* pin wl_1_19
* pin wl_0_19
* pin wl_0_20
* pin wl_1_20
* pin wl_1_21
* pin wl_0_21
* pin wl_0_22
* pin wl_1_22
* pin wl_1_23
* pin wl_0_23
* pin wl_0_24
* pin wl_1_24
* pin wl_1_25
* pin wl_0_25
* pin wl_0_26
* pin wl_1_26
* pin wl_1_27
* pin wl_0_27
* pin wl_0_28
* pin wl_1_28
* pin wl_1_29
* pin wl_0_29
* pin wl_0_30
* pin wl_1_30
* pin wl_1_31
* pin wl_0_31
* pin wl_0_32
* pin wl_1_32
* pin wl_0_33
* pin wl_1_33
* pin wl_0_34
* pin wl_1_34
* pin wl_1_35
* pin wl_0_35
* pin wl_0_36
* pin wl_1_36
* pin wl_1_37
* pin wl_0_37
* pin wl_0_38
* pin wl_1_38
* pin wl_1_39
* pin wl_0_39
* pin wl_0_40
* pin wl_1_40
* pin wl_0_41
* pin wl_1_41
* pin wl_0_42
* pin wl_1_42
* pin wl_0_43
* pin wl_1_43
* pin wl_1_44
* pin wl_0_44
* pin wl_0_45
* pin wl_1_45
* pin wl_0_46
* pin wl_1_46
* pin wl_1_47
* pin wl_0_47
* pin wl_0_48
* pin wl_1_48
* pin wl_1_49
* pin wl_0_49
* pin wl_0_50
* pin wl_1_50
* pin wl_0_51
* pin wl_1_51
* pin wl_0_52
* pin wl_1_52
* pin wl_0_53
* pin wl_1_53
* pin wl_1_54
* pin wl_0_54
* pin wl_1_55
* pin wl_0_55
* pin wl_0_56
* pin wl_1_56
* pin wl_1_57
* pin wl_0_57
* pin wl_0_58
* pin wl_1_58
* pin wl_1_59
* pin wl_0_59
* pin wl_0_60
* pin wl_1_60
* pin wl_1_61
* pin wl_0_61
* pin wl_0_62
* pin wl_1_62
* pin wl_1_63
* pin wl_0_63
* pin rbl_wl_1_0
* pin rbl_wl_1_1
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_replica_bitcell_array_1 1 2 3 4 5 6 7
+ 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33
+ 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59
+ 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85
+ 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108
+ 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127
+ 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146
+ 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165
+ 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184
+ 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266
* net 1 rbl_wl_0_1
* net 2 rbl_wl_0_0
* net 3 bl_0_0
* net 4 bl_1_0
* net 5 br_1_0
* net 6 br_0_0
* net 7 bl_0_1
* net 8 bl_1_1
* net 9 br_1_1
* net 10 br_0_1
* net 11 bl_0_2
* net 12 bl_1_2
* net 13 br_1_2
* net 14 br_0_2
* net 15 bl_0_3
* net 16 bl_1_3
* net 17 br_1_3
* net 18 br_0_3
* net 19 bl_0_4
* net 20 bl_1_4
* net 21 br_1_4
* net 22 br_0_4
* net 23 bl_0_5
* net 24 bl_1_5
* net 25 br_1_5
* net 26 br_0_5
* net 27 bl_0_6
* net 28 bl_1_6
* net 29 br_1_6
* net 30 br_0_6
* net 31 bl_0_7
* net 32 bl_1_7
* net 33 br_1_7
* net 34 br_0_7
* net 35 bl_0_8
* net 36 bl_1_8
* net 37 br_1_8
* net 38 br_0_8
* net 39 bl_0_9
* net 40 bl_1_9
* net 41 br_1_9
* net 42 br_0_9
* net 43 bl_0_10
* net 44 bl_1_10
* net 45 br_1_10
* net 46 br_0_10
* net 47 bl_0_11
* net 48 bl_1_11
* net 49 br_1_11
* net 50 br_0_11
* net 51 bl_0_12
* net 52 bl_1_12
* net 53 br_1_12
* net 54 br_0_12
* net 55 bl_0_13
* net 56 bl_1_13
* net 57 br_1_13
* net 58 br_0_13
* net 59 bl_0_14
* net 60 bl_1_14
* net 61 br_1_14
* net 62 br_0_14
* net 63 bl_0_15
* net 64 bl_1_15
* net 65 br_1_15
* net 66 br_0_15
* net 67 bl_0_16
* net 68 bl_1_16
* net 69 br_1_16
* net 70 br_0_16
* net 71 bl_0_17
* net 72 bl_1_17
* net 73 br_1_17
* net 74 br_0_17
* net 75 bl_0_18
* net 76 bl_1_18
* net 77 br_1_18
* net 78 br_0_18
* net 79 bl_0_19
* net 80 bl_1_19
* net 81 br_1_19
* net 82 br_0_19
* net 83 bl_0_20
* net 84 bl_1_20
* net 85 br_1_20
* net 86 br_0_20
* net 87 bl_0_21
* net 88 bl_1_21
* net 89 br_1_21
* net 90 br_0_21
* net 91 bl_0_22
* net 92 bl_1_22
* net 93 br_1_22
* net 94 br_0_22
* net 95 bl_0_23
* net 96 bl_1_23
* net 97 br_1_23
* net 98 br_0_23
* net 99 bl_0_24
* net 100 bl_1_24
* net 101 br_1_24
* net 102 br_0_24
* net 103 bl_0_25
* net 104 bl_1_25
* net 105 br_1_25
* net 106 br_0_25
* net 107 bl_0_26
* net 108 bl_1_26
* net 109 br_1_26
* net 110 br_0_26
* net 111 bl_0_27
* net 112 bl_1_27
* net 113 br_1_27
* net 114 br_0_27
* net 115 bl_0_28
* net 116 bl_1_28
* net 117 br_1_28
* net 118 br_0_28
* net 119 bl_0_29
* net 120 bl_1_29
* net 121 br_1_29
* net 122 br_0_29
* net 123 bl_0_30
* net 124 bl_1_30
* net 125 br_1_30
* net 126 br_0_30
* net 127 bl_0_31
* net 128 bl_1_31
* net 129 br_1_31
* net 130 br_0_31
* net 131 rbl_bl_0_1
* net 132 rbl_bl_1_1
* net 133 rbl_br_1_1
* net 134 rbl_br_0_1
* net 135 wl_0_0
* net 136 wl_1_0
* net 137 wl_1_1
* net 138 wl_0_1
* net 139 wl_1_2
* net 140 wl_0_2
* net 141 wl_1_3
* net 142 wl_0_3
* net 143 wl_1_4
* net 144 wl_0_4
* net 145 wl_1_5
* net 146 wl_0_5
* net 147 wl_0_6
* net 148 wl_1_6
* net 149 wl_1_7
* net 150 wl_0_7
* net 151 wl_0_8
* net 152 wl_1_8
* net 153 wl_1_9
* net 154 wl_0_9
* net 155 wl_1_10
* net 156 wl_0_10
* net 157 wl_1_11
* net 158 wl_0_11
* net 159 wl_1_12
* net 160 wl_0_12
* net 161 wl_1_13
* net 162 wl_0_13
* net 163 wl_0_14
* net 164 wl_1_14
* net 165 wl_1_15
* net 166 wl_0_15
* net 167 wl_0_16
* net 168 wl_1_16
* net 169 wl_1_17
* net 170 wl_0_17
* net 171 wl_0_18
* net 172 wl_1_18
* net 173 wl_1_19
* net 174 wl_0_19
* net 175 wl_0_20
* net 176 wl_1_20
* net 177 wl_1_21
* net 178 wl_0_21
* net 179 wl_0_22
* net 180 wl_1_22
* net 181 wl_1_23
* net 182 wl_0_23
* net 183 wl_0_24
* net 184 wl_1_24
* net 185 wl_1_25
* net 186 wl_0_25
* net 187 wl_0_26
* net 188 wl_1_26
* net 189 wl_1_27
* net 190 wl_0_27
* net 191 wl_0_28
* net 192 wl_1_28
* net 193 wl_1_29
* net 194 wl_0_29
* net 195 wl_0_30
* net 196 wl_1_30
* net 197 wl_1_31
* net 198 wl_0_31
* net 199 wl_0_32
* net 200 wl_1_32
* net 201 wl_0_33
* net 202 wl_1_33
* net 203 wl_0_34
* net 204 wl_1_34
* net 205 wl_1_35
* net 206 wl_0_35
* net 207 wl_0_36
* net 208 wl_1_36
* net 209 wl_1_37
* net 210 wl_0_37
* net 211 wl_0_38
* net 212 wl_1_38
* net 213 wl_1_39
* net 214 wl_0_39
* net 215 wl_0_40
* net 216 wl_1_40
* net 217 wl_0_41
* net 218 wl_1_41
* net 219 wl_0_42
* net 220 wl_1_42
* net 221 wl_0_43
* net 222 wl_1_43
* net 223 wl_1_44
* net 224 wl_0_44
* net 225 wl_0_45
* net 226 wl_1_45
* net 227 wl_0_46
* net 228 wl_1_46
* net 229 wl_1_47
* net 230 wl_0_47
* net 231 wl_0_48
* net 232 wl_1_48
* net 233 wl_1_49
* net 234 wl_0_49
* net 235 wl_0_50
* net 236 wl_1_50
* net 237 wl_0_51
* net 238 wl_1_51
* net 239 wl_0_52
* net 240 wl_1_52
* net 241 wl_0_53
* net 242 wl_1_53
* net 243 wl_1_54
* net 244 wl_0_54
* net 245 wl_1_55
* net 246 wl_0_55
* net 247 wl_0_56
* net 248 wl_1_56
* net 249 wl_1_57
* net 250 wl_0_57
* net 251 wl_0_58
* net 252 wl_1_58
* net 253 wl_1_59
* net 254 wl_0_59
* net 255 wl_0_60
* net 256 wl_1_60
* net 257 wl_1_61
* net 258 wl_0_61
* net 259 wl_0_62
* net 260 wl_1_62
* net 261 wl_1_63
* net 262 wl_0_63
* net 263 rbl_wl_1_0
* net 264 rbl_wl_1_1
* net 265 vdd
* net 266 gnd
* cell instance $1 r0 *1 37.6,0
X$1 2 1 136 135 138 137 139 140 142 141 143 144 146 145 148 147 150 149 152 151
+ 154 153 155 156 158 157 159 160 162 161 164 163 166 165 168 167 170 169 172
+ 171 174 173 176 175 178 177 180 179 182 181 184 183 186 185 188 187 190 189
+ 192 191 194 193 196 195 131 132 198 197 133 134 200 199 201 202 204 203 206
+ 205 208 207 210 209 212 211 214 213 216 215 217 218 220 219 221 222 223 224
+ 225 226 228 227 230 229 232 231 234 233 236 235 237 238 240 239 241 242 243
+ 244 246 245 248 247 250 249 252 251 254 253 256 255 258 257 260 259 262 261
+ 264 263 265 266 custom_sram_1r1w_32_256_freepdk45_replica_column_0
* cell instance $2 m0 *1 0,1.495
X$2 2 1 265 266 custom_sram_1r1w_32_256_freepdk45_dummy_array_4
* cell instance $3 r0 *1 0,1.495
X$3 140 139 138 137 135 136 143 146 145 144 141 142 149 150 151 152 148 147 156
+ 155 157 158 154 153 163 161 159 164 162 160 168 170 167 169 165 166 176 175
+ 171 174 173 172 179 180 181 182 178 177 186 187 188 183 184 185 191 192 194
+ 190 189 193 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52
+ 53 54 55 56 57 58 59 60 61 62 63 64 65 66 198 197 196 195 67 68 69 70 71 72
+ 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98
+ 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117
+ 118 119 120 121 122 123 124 125 126 127 128 129 130 206 203 202 208 201 205
+ 200 207 199 204 209 214 213 212 210 211 219 220 217 218 215 216 224 223 221
+ 226 222 225 229 230 227 228 231 232 238 237 235 236 233 234 242 244 243 241
+ 240 239 248 245 247 246 250 249 252 256 251 255 254 253 261 262 257 259 260
+ 258 265 266 custom_sram_1r1w_32_256_freepdk45_bitcell_array_0
* cell instance $4 r0 *1 0,97.175
X$4 263 264 265 266 custom_sram_1r1w_32_256_freepdk45_dummy_array_4
.ENDS custom_sram_1r1w_32_256_freepdk45_replica_bitcell_array_1

* cell custom_sram_1r1w_32_256_freepdk45_dummy_array_7
* pin wl_1_0
* pin wl_0_0
* pin wl_0_1
* pin wl_1_1
* pin wl_1_2
* pin wl_0_2
* pin wl_0_3
* pin wl_1_3
* pin wl_1_4
* pin wl_0_4
* pin wl_0_5
* pin wl_1_5
* pin wl_1_6
* pin wl_0_6
* pin wl_0_7
* pin wl_1_7
* pin wl_1_8
* pin wl_0_8
* pin wl_0_9
* pin wl_1_9
* pin wl_1_10
* pin wl_0_10
* pin wl_0_11
* pin wl_1_11
* pin wl_1_12
* pin wl_0_12
* pin wl_0_13
* pin wl_1_13
* pin wl_1_14
* pin wl_0_14
* pin wl_0_15
* pin wl_1_15
* pin wl_1_16
* pin wl_0_16
* pin wl_0_17
* pin wl_1_17
* pin wl_1_18
* pin wl_0_18
* pin wl_0_19
* pin wl_1_19
* pin wl_1_20
* pin wl_0_20
* pin wl_0_21
* pin wl_1_21
* pin wl_1_22
* pin wl_0_22
* pin wl_0_23
* pin wl_1_23
* pin wl_1_24
* pin wl_0_24
* pin wl_0_25
* pin wl_1_25
* pin wl_1_26
* pin wl_0_26
* pin wl_0_27
* pin wl_1_27
* pin wl_1_28
* pin wl_0_28
* pin wl_0_29
* pin wl_1_29
* pin wl_1_30
* pin wl_0_30
* pin wl_0_31
* pin wl_1_31
* pin wl_1_32
* pin wl_0_32
* pin wl_0_33
* pin wl_1_33
* pin wl_1_34
* pin wl_0_34
* pin wl_0_35
* pin wl_1_35
* pin wl_1_36
* pin wl_0_36
* pin wl_0_37
* pin wl_1_37
* pin wl_1_38
* pin wl_0_38
* pin wl_0_39
* pin wl_1_39
* pin wl_1_40
* pin wl_0_40
* pin wl_0_41
* pin wl_1_41
* pin wl_1_42
* pin wl_0_42
* pin wl_0_43
* pin wl_1_43
* pin wl_1_44
* pin wl_0_44
* pin wl_0_45
* pin wl_1_45
* pin wl_1_46
* pin wl_0_46
* pin wl_0_47
* pin wl_1_47
* pin wl_1_48
* pin wl_0_48
* pin wl_0_49
* pin wl_1_49
* pin wl_1_50
* pin wl_0_50
* pin wl_0_51
* pin wl_1_51
* pin wl_1_52
* pin wl_0_52
* pin wl_0_53
* pin wl_1_53
* pin wl_1_54
* pin wl_0_54
* pin wl_0_55
* pin wl_1_55
* pin wl_1_56
* pin wl_0_56
* pin wl_0_57
* pin wl_1_57
* pin wl_1_58
* pin wl_0_58
* pin wl_0_59
* pin wl_1_59
* pin wl_1_60
* pin wl_0_60
* pin wl_0_61
* pin wl_1_61
* pin wl_1_62
* pin wl_0_62
* pin wl_0_63
* pin wl_1_63
* pin wl_1_64
* pin wl_0_64
* pin wl_0_65
* pin wl_1_65
* pin wl_1_66
* pin wl_0_66
* pin wl_0_67
* pin wl_1_67
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_dummy_array_7 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37
+ 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89
+ 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111
+ 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130
+ 131 132 133 134 135 136 137 138
* net 1 wl_1_0
* net 2 wl_0_0
* net 3 wl_0_1
* net 4 wl_1_1
* net 5 wl_1_2
* net 6 wl_0_2
* net 7 wl_0_3
* net 8 wl_1_3
* net 9 wl_1_4
* net 10 wl_0_4
* net 11 wl_0_5
* net 12 wl_1_5
* net 13 wl_1_6
* net 14 wl_0_6
* net 15 wl_0_7
* net 16 wl_1_7
* net 17 wl_1_8
* net 18 wl_0_8
* net 19 wl_0_9
* net 20 wl_1_9
* net 21 wl_1_10
* net 22 wl_0_10
* net 23 wl_0_11
* net 24 wl_1_11
* net 25 wl_1_12
* net 26 wl_0_12
* net 27 wl_0_13
* net 28 wl_1_13
* net 29 wl_1_14
* net 30 wl_0_14
* net 31 wl_0_15
* net 32 wl_1_15
* net 33 wl_1_16
* net 34 wl_0_16
* net 35 wl_0_17
* net 36 wl_1_17
* net 37 wl_1_18
* net 38 wl_0_18
* net 39 wl_0_19
* net 40 wl_1_19
* net 41 wl_1_20
* net 42 wl_0_20
* net 43 wl_0_21
* net 44 wl_1_21
* net 45 wl_1_22
* net 46 wl_0_22
* net 47 wl_0_23
* net 48 wl_1_23
* net 49 wl_1_24
* net 50 wl_0_24
* net 51 wl_0_25
* net 52 wl_1_25
* net 53 wl_1_26
* net 54 wl_0_26
* net 55 wl_0_27
* net 56 wl_1_27
* net 57 wl_1_28
* net 58 wl_0_28
* net 59 wl_0_29
* net 60 wl_1_29
* net 61 wl_1_30
* net 62 wl_0_30
* net 63 wl_0_31
* net 64 wl_1_31
* net 65 wl_1_32
* net 66 wl_0_32
* net 67 wl_0_33
* net 68 wl_1_33
* net 69 wl_1_34
* net 70 wl_0_34
* net 71 wl_0_35
* net 72 wl_1_35
* net 73 wl_1_36
* net 74 wl_0_36
* net 75 wl_0_37
* net 76 wl_1_37
* net 77 wl_1_38
* net 78 wl_0_38
* net 79 wl_0_39
* net 80 wl_1_39
* net 81 wl_1_40
* net 82 wl_0_40
* net 83 wl_0_41
* net 84 wl_1_41
* net 85 wl_1_42
* net 86 wl_0_42
* net 87 wl_0_43
* net 88 wl_1_43
* net 89 wl_1_44
* net 90 wl_0_44
* net 91 wl_0_45
* net 92 wl_1_45
* net 93 wl_1_46
* net 94 wl_0_46
* net 95 wl_0_47
* net 96 wl_1_47
* net 97 wl_1_48
* net 98 wl_0_48
* net 99 wl_0_49
* net 100 wl_1_49
* net 101 wl_1_50
* net 102 wl_0_50
* net 103 wl_0_51
* net 104 wl_1_51
* net 105 wl_1_52
* net 106 wl_0_52
* net 107 wl_0_53
* net 108 wl_1_53
* net 109 wl_1_54
* net 110 wl_0_54
* net 111 wl_0_55
* net 112 wl_1_55
* net 113 wl_1_56
* net 114 wl_0_56
* net 115 wl_0_57
* net 116 wl_1_57
* net 117 wl_1_58
* net 118 wl_0_58
* net 119 wl_0_59
* net 120 wl_1_59
* net 121 wl_1_60
* net 122 wl_0_60
* net 123 wl_0_61
* net 124 wl_1_61
* net 125 wl_1_62
* net 126 wl_0_62
* net 127 wl_0_63
* net 128 wl_1_63
* net 129 wl_1_64
* net 130 wl_0_64
* net 131 wl_0_65
* net 132 wl_1_65
* net 133 wl_1_66
* net 134 wl_0_66
* net 135 wl_0_67
* net 136 wl_1_67
* net 137 vdd
* net 138 gnd
* cell instance $1 r0 *1 0,0
X$1 1 2 137 138 dummy_cell_2rw
* cell instance $2 m0 *1 0,2.99
X$2 4 3 137 138 dummy_cell_2rw
* cell instance $3 r0 *1 0,2.99
X$3 5 6 137 138 dummy_cell_2rw
* cell instance $4 m0 *1 0,5.98
X$4 8 7 137 138 dummy_cell_2rw
* cell instance $5 r0 *1 0,5.98
X$5 9 10 137 138 dummy_cell_2rw
* cell instance $6 m0 *1 0,8.97
X$6 12 11 137 138 dummy_cell_2rw
* cell instance $7 r0 *1 0,8.97
X$7 13 14 137 138 dummy_cell_2rw
* cell instance $8 m0 *1 0,11.96
X$8 16 15 137 138 dummy_cell_2rw
* cell instance $9 r0 *1 0,11.96
X$9 17 18 137 138 dummy_cell_2rw
* cell instance $10 m0 *1 0,14.95
X$10 20 19 137 138 dummy_cell_2rw
* cell instance $11 r0 *1 0,14.95
X$11 21 22 137 138 dummy_cell_2rw
* cell instance $12 m0 *1 0,17.94
X$12 24 23 137 138 dummy_cell_2rw
* cell instance $13 r0 *1 0,17.94
X$13 25 26 137 138 dummy_cell_2rw
* cell instance $14 m0 *1 0,20.93
X$14 28 27 137 138 dummy_cell_2rw
* cell instance $15 r0 *1 0,20.93
X$15 29 30 137 138 dummy_cell_2rw
* cell instance $16 m0 *1 0,23.92
X$16 32 31 137 138 dummy_cell_2rw
* cell instance $17 r0 *1 0,23.92
X$17 33 34 137 138 dummy_cell_2rw
* cell instance $18 m0 *1 0,26.91
X$18 36 35 137 138 dummy_cell_2rw
* cell instance $19 r0 *1 0,26.91
X$19 37 38 137 138 dummy_cell_2rw
* cell instance $20 m0 *1 0,29.9
X$20 40 39 137 138 dummy_cell_2rw
* cell instance $21 r0 *1 0,29.9
X$21 41 42 137 138 dummy_cell_2rw
* cell instance $22 m0 *1 0,32.89
X$22 44 43 137 138 dummy_cell_2rw
* cell instance $23 r0 *1 0,32.89
X$23 45 46 137 138 dummy_cell_2rw
* cell instance $24 m0 *1 0,35.88
X$24 48 47 137 138 dummy_cell_2rw
* cell instance $25 r0 *1 0,35.88
X$25 49 50 137 138 dummy_cell_2rw
* cell instance $26 m0 *1 0,38.87
X$26 52 51 137 138 dummy_cell_2rw
* cell instance $27 r0 *1 0,38.87
X$27 53 54 137 138 dummy_cell_2rw
* cell instance $28 m0 *1 0,41.86
X$28 56 55 137 138 dummy_cell_2rw
* cell instance $29 r0 *1 0,41.86
X$29 57 58 137 138 dummy_cell_2rw
* cell instance $30 m0 *1 0,44.85
X$30 60 59 137 138 dummy_cell_2rw
* cell instance $31 r0 *1 0,44.85
X$31 61 62 137 138 dummy_cell_2rw
* cell instance $32 m0 *1 0,47.84
X$32 64 63 137 138 dummy_cell_2rw
* cell instance $33 r0 *1 0,47.84
X$33 65 66 137 138 dummy_cell_2rw
* cell instance $34 m0 *1 0,50.83
X$34 68 67 137 138 dummy_cell_2rw
* cell instance $35 r0 *1 0,50.83
X$35 69 70 137 138 dummy_cell_2rw
* cell instance $36 m0 *1 0,53.82
X$36 72 71 137 138 dummy_cell_2rw
* cell instance $37 r0 *1 0,53.82
X$37 73 74 137 138 dummy_cell_2rw
* cell instance $38 m0 *1 0,56.81
X$38 76 75 137 138 dummy_cell_2rw
* cell instance $39 r0 *1 0,56.81
X$39 77 78 137 138 dummy_cell_2rw
* cell instance $40 m0 *1 0,59.8
X$40 80 79 137 138 dummy_cell_2rw
* cell instance $41 r0 *1 0,59.8
X$41 81 82 137 138 dummy_cell_2rw
* cell instance $42 m0 *1 0,62.79
X$42 84 83 137 138 dummy_cell_2rw
* cell instance $43 r0 *1 0,62.79
X$43 85 86 137 138 dummy_cell_2rw
* cell instance $44 m0 *1 0,65.78
X$44 88 87 137 138 dummy_cell_2rw
* cell instance $45 r0 *1 0,65.78
X$45 89 90 137 138 dummy_cell_2rw
* cell instance $46 m0 *1 0,68.77
X$46 92 91 137 138 dummy_cell_2rw
* cell instance $47 r0 *1 0,68.77
X$47 93 94 137 138 dummy_cell_2rw
* cell instance $48 m0 *1 0,71.76
X$48 96 95 137 138 dummy_cell_2rw
* cell instance $49 r0 *1 0,71.76
X$49 97 98 137 138 dummy_cell_2rw
* cell instance $50 m0 *1 0,74.75
X$50 100 99 137 138 dummy_cell_2rw
* cell instance $51 r0 *1 0,74.75
X$51 101 102 137 138 dummy_cell_2rw
* cell instance $52 m0 *1 0,77.74
X$52 104 103 137 138 dummy_cell_2rw
* cell instance $53 r0 *1 0,77.74
X$53 105 106 137 138 dummy_cell_2rw
* cell instance $54 m0 *1 0,80.73
X$54 108 107 137 138 dummy_cell_2rw
* cell instance $55 r0 *1 0,80.73
X$55 109 110 137 138 dummy_cell_2rw
* cell instance $56 m0 *1 0,83.72
X$56 112 111 137 138 dummy_cell_2rw
* cell instance $57 r0 *1 0,83.72
X$57 113 114 137 138 dummy_cell_2rw
* cell instance $58 m0 *1 0,86.71
X$58 116 115 137 138 dummy_cell_2rw
* cell instance $59 r0 *1 0,86.71
X$59 117 118 137 138 dummy_cell_2rw
* cell instance $60 m0 *1 0,89.7
X$60 120 119 137 138 dummy_cell_2rw
* cell instance $61 r0 *1 0,89.7
X$61 121 122 137 138 dummy_cell_2rw
* cell instance $62 m0 *1 0,92.69
X$62 124 123 137 138 dummy_cell_2rw
* cell instance $63 r0 *1 0,92.69
X$63 125 126 137 138 dummy_cell_2rw
* cell instance $64 m0 *1 0,95.68
X$64 128 127 137 138 dummy_cell_2rw
* cell instance $65 r0 *1 0,95.68
X$65 129 130 137 138 dummy_cell_2rw
* cell instance $66 m0 *1 0,98.67
X$66 132 131 137 138 dummy_cell_2rw
* cell instance $67 r0 *1 0,98.67
X$67 133 134 137 138 dummy_cell_2rw
* cell instance $68 m0 *1 0,101.66
X$68 136 135 137 138 dummy_cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_dummy_array_7

* cell custom_sram_1r1w_32_256_freepdk45_dummy_array_5
* pin wl_0_0
* pin wl_1_0
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_dummy_array_5 1 2 3 4
* net 1 wl_0_0
* net 2 wl_1_0
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 dummy_cell_2rw
* cell instance $2 r0 *1 1.175,0
X$2 2 1 3 4 dummy_cell_2rw
* cell instance $3 r0 *1 2.35,0
X$3 2 1 3 4 dummy_cell_2rw
* cell instance $4 r0 *1 3.525,0
X$4 2 1 3 4 dummy_cell_2rw
* cell instance $5 r0 *1 4.7,0
X$5 2 1 3 4 dummy_cell_2rw
* cell instance $6 r0 *1 5.875,0
X$6 2 1 3 4 dummy_cell_2rw
* cell instance $7 r0 *1 7.05,0
X$7 2 1 3 4 dummy_cell_2rw
* cell instance $8 r0 *1 8.225,0
X$8 2 1 3 4 dummy_cell_2rw
* cell instance $9 r0 *1 9.4,0
X$9 2 1 3 4 dummy_cell_2rw
* cell instance $10 r0 *1 10.575,0
X$10 2 1 3 4 dummy_cell_2rw
* cell instance $11 r0 *1 11.75,0
X$11 2 1 3 4 dummy_cell_2rw
* cell instance $12 r0 *1 12.925,0
X$12 2 1 3 4 dummy_cell_2rw
* cell instance $13 r0 *1 14.1,0
X$13 2 1 3 4 dummy_cell_2rw
* cell instance $14 r0 *1 15.275,0
X$14 2 1 3 4 dummy_cell_2rw
* cell instance $15 r0 *1 16.45,0
X$15 2 1 3 4 dummy_cell_2rw
* cell instance $16 r0 *1 17.625,0
X$16 2 1 3 4 dummy_cell_2rw
* cell instance $17 r0 *1 18.8,0
X$17 2 1 3 4 dummy_cell_2rw
* cell instance $18 r0 *1 19.975,0
X$18 2 1 3 4 dummy_cell_2rw
* cell instance $19 r0 *1 21.15,0
X$19 2 1 3 4 dummy_cell_2rw
* cell instance $20 r0 *1 22.325,0
X$20 2 1 3 4 dummy_cell_2rw
* cell instance $21 r0 *1 23.5,0
X$21 2 1 3 4 dummy_cell_2rw
* cell instance $22 r0 *1 24.675,0
X$22 2 1 3 4 dummy_cell_2rw
* cell instance $23 r0 *1 25.85,0
X$23 2 1 3 4 dummy_cell_2rw
* cell instance $24 r0 *1 27.025,0
X$24 2 1 3 4 dummy_cell_2rw
* cell instance $25 r0 *1 28.2,0
X$25 2 1 3 4 dummy_cell_2rw
* cell instance $26 r0 *1 29.375,0
X$26 2 1 3 4 dummy_cell_2rw
* cell instance $27 r0 *1 30.55,0
X$27 2 1 3 4 dummy_cell_2rw
* cell instance $28 r0 *1 31.725,0
X$28 2 1 3 4 dummy_cell_2rw
* cell instance $29 r0 *1 32.9,0
X$29 2 1 3 4 dummy_cell_2rw
* cell instance $30 r0 *1 34.075,0
X$30 2 1 3 4 dummy_cell_2rw
* cell instance $31 r0 *1 35.25,0
X$31 2 1 3 4 dummy_cell_2rw
* cell instance $32 r0 *1 36.425,0
X$32 2 1 3 4 dummy_cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_dummy_array_5

* cell custom_sram_1r1w_32_256_freepdk45_dummy_array_6
* pin wl_0_0
* pin wl_1_0
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_dummy_array_6 1 2 3 4
* net 1 wl_0_0
* net 2 wl_1_0
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 dummy_cell_2rw
* cell instance $2 r0 *1 1.175,0
X$2 2 1 3 4 dummy_cell_2rw
* cell instance $3 r0 *1 2.35,0
X$3 2 1 3 4 dummy_cell_2rw
* cell instance $4 r0 *1 3.525,0
X$4 2 1 3 4 dummy_cell_2rw
* cell instance $5 r0 *1 4.7,0
X$5 2 1 3 4 dummy_cell_2rw
* cell instance $6 r0 *1 5.875,0
X$6 2 1 3 4 dummy_cell_2rw
* cell instance $7 r0 *1 7.05,0
X$7 2 1 3 4 dummy_cell_2rw
* cell instance $8 r0 *1 8.225,0
X$8 2 1 3 4 dummy_cell_2rw
* cell instance $9 r0 *1 9.4,0
X$9 2 1 3 4 dummy_cell_2rw
* cell instance $10 r0 *1 10.575,0
X$10 2 1 3 4 dummy_cell_2rw
* cell instance $11 r0 *1 11.75,0
X$11 2 1 3 4 dummy_cell_2rw
* cell instance $12 r0 *1 12.925,0
X$12 2 1 3 4 dummy_cell_2rw
* cell instance $13 r0 *1 14.1,0
X$13 2 1 3 4 dummy_cell_2rw
* cell instance $14 r0 *1 15.275,0
X$14 2 1 3 4 dummy_cell_2rw
* cell instance $15 r0 *1 16.45,0
X$15 2 1 3 4 dummy_cell_2rw
* cell instance $16 r0 *1 17.625,0
X$16 2 1 3 4 dummy_cell_2rw
* cell instance $17 r0 *1 18.8,0
X$17 2 1 3 4 dummy_cell_2rw
* cell instance $18 r0 *1 19.975,0
X$18 2 1 3 4 dummy_cell_2rw
* cell instance $19 r0 *1 21.15,0
X$19 2 1 3 4 dummy_cell_2rw
* cell instance $20 r0 *1 22.325,0
X$20 2 1 3 4 dummy_cell_2rw
* cell instance $21 r0 *1 23.5,0
X$21 2 1 3 4 dummy_cell_2rw
* cell instance $22 r0 *1 24.675,0
X$22 2 1 3 4 dummy_cell_2rw
* cell instance $23 r0 *1 25.85,0
X$23 2 1 3 4 dummy_cell_2rw
* cell instance $24 r0 *1 27.025,0
X$24 2 1 3 4 dummy_cell_2rw
* cell instance $25 r0 *1 28.2,0
X$25 2 1 3 4 dummy_cell_2rw
* cell instance $26 r0 *1 29.375,0
X$26 2 1 3 4 dummy_cell_2rw
* cell instance $27 r0 *1 30.55,0
X$27 2 1 3 4 dummy_cell_2rw
* cell instance $28 r0 *1 31.725,0
X$28 2 1 3 4 dummy_cell_2rw
* cell instance $29 r0 *1 32.9,0
X$29 2 1 3 4 dummy_cell_2rw
* cell instance $30 r0 *1 34.075,0
X$30 2 1 3 4 dummy_cell_2rw
* cell instance $31 r0 *1 35.25,0
X$31 2 1 3 4 dummy_cell_2rw
* cell instance $32 r0 *1 36.425,0
X$32 2 1 3 4 dummy_cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_dummy_array_6

* cell custom_sram_1r1w_32_256_freepdk45_replica_bitcell_array_0
* pin rbl_wl_0_0
* pin rbl_wl_0_1
* pin bl_0_0
* pin bl_1_0
* pin br_1_0
* pin br_0_0
* pin bl_0_1
* pin bl_1_1
* pin br_1_1
* pin br_0_1
* pin bl_0_2
* pin bl_1_2
* pin br_1_2
* pin br_0_2
* pin bl_0_3
* pin bl_1_3
* pin br_1_3
* pin br_0_3
* pin bl_0_4
* pin bl_1_4
* pin br_1_4
* pin br_0_4
* pin bl_0_5
* pin bl_1_5
* pin br_1_5
* pin br_0_5
* pin bl_0_6
* pin bl_1_6
* pin br_1_6
* pin br_0_6
* pin bl_0_7
* pin bl_1_7
* pin br_1_7
* pin br_0_7
* pin bl_0_8
* pin bl_1_8
* pin br_1_8
* pin br_0_8
* pin bl_0_9
* pin bl_1_9
* pin br_1_9
* pin br_0_9
* pin bl_0_10
* pin bl_1_10
* pin br_1_10
* pin br_0_10
* pin bl_0_11
* pin bl_1_11
* pin br_1_11
* pin br_0_11
* pin bl_0_12
* pin bl_1_12
* pin br_1_12
* pin br_0_12
* pin bl_0_13
* pin bl_1_13
* pin br_1_13
* pin br_0_13
* pin bl_0_14
* pin bl_1_14
* pin br_1_14
* pin br_0_14
* pin bl_0_15
* pin bl_1_15
* pin br_1_15
* pin br_0_15
* pin bl_0_16
* pin bl_1_16
* pin br_1_16
* pin br_0_16
* pin bl_0_17
* pin bl_1_17
* pin br_1_17
* pin br_0_17
* pin bl_0_18
* pin bl_1_18
* pin br_1_18
* pin br_0_18
* pin bl_0_19
* pin bl_1_19
* pin br_1_19
* pin br_0_19
* pin bl_0_20
* pin bl_1_20
* pin br_1_20
* pin br_0_20
* pin bl_0_21
* pin bl_1_21
* pin br_1_21
* pin br_0_21
* pin bl_0_22
* pin bl_1_22
* pin br_1_22
* pin br_0_22
* pin bl_0_23
* pin bl_1_23
* pin br_1_23
* pin br_0_23
* pin bl_0_24
* pin bl_1_24
* pin br_1_24
* pin br_0_24
* pin bl_0_25
* pin bl_1_25
* pin br_1_25
* pin br_0_25
* pin bl_0_26
* pin bl_1_26
* pin br_1_26
* pin br_0_26
* pin bl_0_27
* pin bl_1_27
* pin br_1_27
* pin br_0_27
* pin bl_0_28
* pin bl_1_28
* pin br_1_28
* pin br_0_28
* pin bl_0_29
* pin bl_1_29
* pin br_1_29
* pin br_0_29
* pin bl_0_30
* pin bl_1_30
* pin br_1_30
* pin br_0_30
* pin bl_0_31
* pin bl_1_31
* pin br_1_31
* pin br_0_31
* pin wl_1_0
* pin wl_0_0
* pin wl_0_1
* pin wl_1_1
* pin wl_0_2
* pin wl_1_2
* pin wl_1_3
* pin wl_0_3
* pin wl_0_4
* pin wl_1_4
* pin wl_1_5
* pin wl_0_5
* pin wl_1_6
* pin wl_0_6
* pin wl_1_7
* pin wl_0_7
* pin wl_1_8
* pin wl_0_8
* pin wl_1_9
* pin wl_0_9
* pin wl_1_10
* pin wl_0_10
* pin wl_0_11
* pin wl_1_11
* pin wl_0_12
* pin wl_1_12
* pin wl_1_13
* pin wl_0_13
* pin wl_0_14
* pin wl_1_14
* pin wl_0_15
* pin wl_1_15
* pin wl_0_16
* pin wl_1_16
* pin wl_1_17
* pin wl_0_17
* pin wl_1_18
* pin wl_0_18
* pin wl_1_19
* pin wl_0_19
* pin wl_1_20
* pin wl_0_20
* pin wl_0_21
* pin wl_1_21
* pin wl_1_22
* pin wl_0_22
* pin wl_0_23
* pin wl_1_23
* pin wl_1_24
* pin wl_0_24
* pin wl_1_25
* pin wl_0_25
* pin wl_0_26
* pin wl_1_26
* pin wl_1_27
* pin wl_0_27
* pin wl_1_28
* pin wl_0_28
* pin wl_1_29
* pin wl_0_29
* pin wl_1_30
* pin wl_0_30
* pin wl_1_31
* pin wl_0_31
* pin wl_1_32
* pin wl_0_32
* pin wl_0_33
* pin wl_1_33
* pin wl_0_34
* pin wl_1_34
* pin wl_1_35
* pin wl_0_35
* pin wl_0_36
* pin wl_1_36
* pin wl_1_37
* pin wl_0_37
* pin wl_0_38
* pin wl_1_38
* pin wl_1_39
* pin wl_0_39
* pin wl_0_40
* pin wl_1_40
* pin wl_1_41
* pin wl_0_41
* pin wl_0_42
* pin wl_1_42
* pin wl_1_43
* pin wl_0_43
* pin wl_1_44
* pin wl_0_44
* pin wl_1_45
* pin wl_0_45
* pin wl_1_46
* pin wl_0_46
* pin wl_1_47
* pin wl_0_47
* pin wl_1_48
* pin wl_0_48
* pin wl_1_49
* pin wl_0_49
* pin wl_0_50
* pin wl_1_50
* pin wl_1_51
* pin wl_0_51
* pin wl_0_52
* pin wl_1_52
* pin wl_0_53
* pin wl_1_53
* pin wl_1_54
* pin wl_0_54
* pin wl_0_55
* pin wl_1_55
* pin wl_0_56
* pin wl_1_56
* pin wl_1_57
* pin wl_0_57
* pin wl_1_58
* pin wl_0_58
* pin wl_1_59
* pin wl_0_59
* pin wl_0_60
* pin wl_1_60
* pin wl_0_61
* pin wl_1_61
* pin wl_1_62
* pin wl_0_62
* pin wl_1_63
* pin wl_0_63
* pin rbl_wl_1_0
* pin rbl_wl_1_1
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_replica_bitcell_array_0 1 2 3 4 5 6 7
+ 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33
+ 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59
+ 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85
+ 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108
+ 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127
+ 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146
+ 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165
+ 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184
+ 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262
* net 1 rbl_wl_0_0
* net 2 rbl_wl_0_1
* net 3 bl_0_0
* net 4 bl_1_0
* net 5 br_1_0
* net 6 br_0_0
* net 7 bl_0_1
* net 8 bl_1_1
* net 9 br_1_1
* net 10 br_0_1
* net 11 bl_0_2
* net 12 bl_1_2
* net 13 br_1_2
* net 14 br_0_2
* net 15 bl_0_3
* net 16 bl_1_3
* net 17 br_1_3
* net 18 br_0_3
* net 19 bl_0_4
* net 20 bl_1_4
* net 21 br_1_4
* net 22 br_0_4
* net 23 bl_0_5
* net 24 bl_1_5
* net 25 br_1_5
* net 26 br_0_5
* net 27 bl_0_6
* net 28 bl_1_6
* net 29 br_1_6
* net 30 br_0_6
* net 31 bl_0_7
* net 32 bl_1_7
* net 33 br_1_7
* net 34 br_0_7
* net 35 bl_0_8
* net 36 bl_1_8
* net 37 br_1_8
* net 38 br_0_8
* net 39 bl_0_9
* net 40 bl_1_9
* net 41 br_1_9
* net 42 br_0_9
* net 43 bl_0_10
* net 44 bl_1_10
* net 45 br_1_10
* net 46 br_0_10
* net 47 bl_0_11
* net 48 bl_1_11
* net 49 br_1_11
* net 50 br_0_11
* net 51 bl_0_12
* net 52 bl_1_12
* net 53 br_1_12
* net 54 br_0_12
* net 55 bl_0_13
* net 56 bl_1_13
* net 57 br_1_13
* net 58 br_0_13
* net 59 bl_0_14
* net 60 bl_1_14
* net 61 br_1_14
* net 62 br_0_14
* net 63 bl_0_15
* net 64 bl_1_15
* net 65 br_1_15
* net 66 br_0_15
* net 67 bl_0_16
* net 68 bl_1_16
* net 69 br_1_16
* net 70 br_0_16
* net 71 bl_0_17
* net 72 bl_1_17
* net 73 br_1_17
* net 74 br_0_17
* net 75 bl_0_18
* net 76 bl_1_18
* net 77 br_1_18
* net 78 br_0_18
* net 79 bl_0_19
* net 80 bl_1_19
* net 81 br_1_19
* net 82 br_0_19
* net 83 bl_0_20
* net 84 bl_1_20
* net 85 br_1_20
* net 86 br_0_20
* net 87 bl_0_21
* net 88 bl_1_21
* net 89 br_1_21
* net 90 br_0_21
* net 91 bl_0_22
* net 92 bl_1_22
* net 93 br_1_22
* net 94 br_0_22
* net 95 bl_0_23
* net 96 bl_1_23
* net 97 br_1_23
* net 98 br_0_23
* net 99 bl_0_24
* net 100 bl_1_24
* net 101 br_1_24
* net 102 br_0_24
* net 103 bl_0_25
* net 104 bl_1_25
* net 105 br_1_25
* net 106 br_0_25
* net 107 bl_0_26
* net 108 bl_1_26
* net 109 br_1_26
* net 110 br_0_26
* net 111 bl_0_27
* net 112 bl_1_27
* net 113 br_1_27
* net 114 br_0_27
* net 115 bl_0_28
* net 116 bl_1_28
* net 117 br_1_28
* net 118 br_0_28
* net 119 bl_0_29
* net 120 bl_1_29
* net 121 br_1_29
* net 122 br_0_29
* net 123 bl_0_30
* net 124 bl_1_30
* net 125 br_1_30
* net 126 br_0_30
* net 127 bl_0_31
* net 128 bl_1_31
* net 129 br_1_31
* net 130 br_0_31
* net 131 wl_1_0
* net 132 wl_0_0
* net 133 wl_0_1
* net 134 wl_1_1
* net 135 wl_0_2
* net 136 wl_1_2
* net 137 wl_1_3
* net 138 wl_0_3
* net 139 wl_0_4
* net 140 wl_1_4
* net 141 wl_1_5
* net 142 wl_0_5
* net 143 wl_1_6
* net 144 wl_0_6
* net 145 wl_1_7
* net 146 wl_0_7
* net 147 wl_1_8
* net 148 wl_0_8
* net 149 wl_1_9
* net 150 wl_0_9
* net 151 wl_1_10
* net 152 wl_0_10
* net 153 wl_0_11
* net 154 wl_1_11
* net 155 wl_0_12
* net 156 wl_1_12
* net 157 wl_1_13
* net 158 wl_0_13
* net 159 wl_0_14
* net 160 wl_1_14
* net 161 wl_0_15
* net 162 wl_1_15
* net 163 wl_0_16
* net 164 wl_1_16
* net 165 wl_1_17
* net 166 wl_0_17
* net 167 wl_1_18
* net 168 wl_0_18
* net 169 wl_1_19
* net 170 wl_0_19
* net 171 wl_1_20
* net 172 wl_0_20
* net 173 wl_0_21
* net 174 wl_1_21
* net 175 wl_1_22
* net 176 wl_0_22
* net 177 wl_0_23
* net 178 wl_1_23
* net 179 wl_1_24
* net 180 wl_0_24
* net 181 wl_1_25
* net 182 wl_0_25
* net 183 wl_0_26
* net 184 wl_1_26
* net 185 wl_1_27
* net 186 wl_0_27
* net 187 wl_1_28
* net 188 wl_0_28
* net 189 wl_1_29
* net 190 wl_0_29
* net 191 wl_1_30
* net 192 wl_0_30
* net 193 wl_1_31
* net 194 wl_0_31
* net 195 wl_1_32
* net 196 wl_0_32
* net 197 wl_0_33
* net 198 wl_1_33
* net 199 wl_0_34
* net 200 wl_1_34
* net 201 wl_1_35
* net 202 wl_0_35
* net 203 wl_0_36
* net 204 wl_1_36
* net 205 wl_1_37
* net 206 wl_0_37
* net 207 wl_0_38
* net 208 wl_1_38
* net 209 wl_1_39
* net 210 wl_0_39
* net 211 wl_0_40
* net 212 wl_1_40
* net 213 wl_1_41
* net 214 wl_0_41
* net 215 wl_0_42
* net 216 wl_1_42
* net 217 wl_1_43
* net 218 wl_0_43
* net 219 wl_1_44
* net 220 wl_0_44
* net 221 wl_1_45
* net 222 wl_0_45
* net 223 wl_1_46
* net 224 wl_0_46
* net 225 wl_1_47
* net 226 wl_0_47
* net 227 wl_1_48
* net 228 wl_0_48
* net 229 wl_1_49
* net 230 wl_0_49
* net 231 wl_0_50
* net 232 wl_1_50
* net 233 wl_1_51
* net 234 wl_0_51
* net 235 wl_0_52
* net 236 wl_1_52
* net 237 wl_0_53
* net 238 wl_1_53
* net 239 wl_1_54
* net 240 wl_0_54
* net 241 wl_0_55
* net 242 wl_1_55
* net 243 wl_0_56
* net 244 wl_1_56
* net 245 wl_1_57
* net 246 wl_0_57
* net 247 wl_1_58
* net 248 wl_0_58
* net 249 wl_1_59
* net 250 wl_0_59
* net 251 wl_0_60
* net 252 wl_1_60
* net 253 wl_0_61
* net 254 wl_1_61
* net 255 wl_1_62
* net 256 wl_0_62
* net 257 wl_1_63
* net 258 wl_0_63
* net 259 rbl_wl_1_0
* net 260 rbl_wl_1_1
* net 261 vdd
* net 262 gnd
* cell instance $1 m0 *1 0,1.495
X$1 1 2 261 262 custom_sram_1r1w_32_256_freepdk45_dummy_array_4
* cell instance $2 r0 *1 0,1.495
X$2 135 136 133 134 132 131 140 142 141 139 137 138 145 146 148 147 143 144 152
+ 151 154 153 150 149 159 157 156 160 158 155 164 166 163 165 162 161 171 172
+ 168 170 169 167 176 175 178 177 173 174 182 183 184 180 179 181 188 187 190
+ 186 185 189 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52
+ 53 54 55 56 57 58 59 60 61 62 63 64 65 66 194 193 191 192 67 68 69 70 71 72
+ 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98
+ 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117
+ 118 119 120 121 122 123 124 125 126 127 128 129 130 202 199 198 204 197 201
+ 195 203 196 200 205 210 209 208 206 207 215 216 214 213 211 212 220 219 218
+ 221 217 222 225 226 224 223 228 227 233 234 231 232 229 230 238 240 239 237
+ 236 235 244 242 243 241 246 245 247 252 248 251 250 249 257 258 254 256 255
+ 253 261 262 custom_sram_1r1w_32_256_freepdk45_bitcell_array_0
* cell instance $3 r0 *1 0,97.175
X$3 259 260 261 262 custom_sram_1r1w_32_256_freepdk45_dummy_array_4
.ENDS custom_sram_1r1w_32_256_freepdk45_replica_bitcell_array_0

* cell custom_sram_1r1w_32_256_freepdk45_dummy_array_3
* pin wl_1_0
* pin wl_0_0
* pin wl_0_1
* pin wl_1_1
* pin wl_1_2
* pin wl_0_2
* pin wl_0_3
* pin wl_1_3
* pin wl_1_4
* pin wl_0_4
* pin wl_0_5
* pin wl_1_5
* pin wl_1_6
* pin wl_0_6
* pin wl_0_7
* pin wl_1_7
* pin wl_1_8
* pin wl_0_8
* pin wl_0_9
* pin wl_1_9
* pin wl_1_10
* pin wl_0_10
* pin wl_0_11
* pin wl_1_11
* pin wl_1_12
* pin wl_0_12
* pin wl_0_13
* pin wl_1_13
* pin wl_1_14
* pin wl_0_14
* pin wl_0_15
* pin wl_1_15
* pin wl_1_16
* pin wl_0_16
* pin wl_0_17
* pin wl_1_17
* pin wl_1_18
* pin wl_0_18
* pin wl_0_19
* pin wl_1_19
* pin wl_1_20
* pin wl_0_20
* pin wl_0_21
* pin wl_1_21
* pin wl_1_22
* pin wl_0_22
* pin wl_0_23
* pin wl_1_23
* pin wl_1_24
* pin wl_0_24
* pin wl_0_25
* pin wl_1_25
* pin wl_1_26
* pin wl_0_26
* pin wl_0_27
* pin wl_1_27
* pin wl_1_28
* pin wl_0_28
* pin wl_0_29
* pin wl_1_29
* pin wl_1_30
* pin wl_0_30
* pin wl_0_31
* pin wl_1_31
* pin wl_1_32
* pin wl_0_32
* pin wl_0_33
* pin wl_1_33
* pin wl_1_34
* pin wl_0_34
* pin wl_0_35
* pin wl_1_35
* pin wl_1_36
* pin wl_0_36
* pin wl_0_37
* pin wl_1_37
* pin wl_1_38
* pin wl_0_38
* pin wl_0_39
* pin wl_1_39
* pin wl_1_40
* pin wl_0_40
* pin wl_0_41
* pin wl_1_41
* pin wl_1_42
* pin wl_0_42
* pin wl_0_43
* pin wl_1_43
* pin wl_1_44
* pin wl_0_44
* pin wl_0_45
* pin wl_1_45
* pin wl_1_46
* pin wl_0_46
* pin wl_0_47
* pin wl_1_47
* pin wl_1_48
* pin wl_0_48
* pin wl_0_49
* pin wl_1_49
* pin wl_1_50
* pin wl_0_50
* pin wl_0_51
* pin wl_1_51
* pin wl_1_52
* pin wl_0_52
* pin wl_0_53
* pin wl_1_53
* pin wl_1_54
* pin wl_0_54
* pin wl_0_55
* pin wl_1_55
* pin wl_1_56
* pin wl_0_56
* pin wl_0_57
* pin wl_1_57
* pin wl_1_58
* pin wl_0_58
* pin wl_0_59
* pin wl_1_59
* pin wl_1_60
* pin wl_0_60
* pin wl_0_61
* pin wl_1_61
* pin wl_1_62
* pin wl_0_62
* pin wl_0_63
* pin wl_1_63
* pin wl_1_64
* pin wl_0_64
* pin wl_0_65
* pin wl_1_65
* pin wl_1_66
* pin wl_0_66
* pin wl_0_67
* pin wl_1_67
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_dummy_array_3 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37
+ 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89
+ 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111
+ 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130
+ 131 132 133 134 135 136 137 138
* net 1 wl_1_0
* net 2 wl_0_0
* net 3 wl_0_1
* net 4 wl_1_1
* net 5 wl_1_2
* net 6 wl_0_2
* net 7 wl_0_3
* net 8 wl_1_3
* net 9 wl_1_4
* net 10 wl_0_4
* net 11 wl_0_5
* net 12 wl_1_5
* net 13 wl_1_6
* net 14 wl_0_6
* net 15 wl_0_7
* net 16 wl_1_7
* net 17 wl_1_8
* net 18 wl_0_8
* net 19 wl_0_9
* net 20 wl_1_9
* net 21 wl_1_10
* net 22 wl_0_10
* net 23 wl_0_11
* net 24 wl_1_11
* net 25 wl_1_12
* net 26 wl_0_12
* net 27 wl_0_13
* net 28 wl_1_13
* net 29 wl_1_14
* net 30 wl_0_14
* net 31 wl_0_15
* net 32 wl_1_15
* net 33 wl_1_16
* net 34 wl_0_16
* net 35 wl_0_17
* net 36 wl_1_17
* net 37 wl_1_18
* net 38 wl_0_18
* net 39 wl_0_19
* net 40 wl_1_19
* net 41 wl_1_20
* net 42 wl_0_20
* net 43 wl_0_21
* net 44 wl_1_21
* net 45 wl_1_22
* net 46 wl_0_22
* net 47 wl_0_23
* net 48 wl_1_23
* net 49 wl_1_24
* net 50 wl_0_24
* net 51 wl_0_25
* net 52 wl_1_25
* net 53 wl_1_26
* net 54 wl_0_26
* net 55 wl_0_27
* net 56 wl_1_27
* net 57 wl_1_28
* net 58 wl_0_28
* net 59 wl_0_29
* net 60 wl_1_29
* net 61 wl_1_30
* net 62 wl_0_30
* net 63 wl_0_31
* net 64 wl_1_31
* net 65 wl_1_32
* net 66 wl_0_32
* net 67 wl_0_33
* net 68 wl_1_33
* net 69 wl_1_34
* net 70 wl_0_34
* net 71 wl_0_35
* net 72 wl_1_35
* net 73 wl_1_36
* net 74 wl_0_36
* net 75 wl_0_37
* net 76 wl_1_37
* net 77 wl_1_38
* net 78 wl_0_38
* net 79 wl_0_39
* net 80 wl_1_39
* net 81 wl_1_40
* net 82 wl_0_40
* net 83 wl_0_41
* net 84 wl_1_41
* net 85 wl_1_42
* net 86 wl_0_42
* net 87 wl_0_43
* net 88 wl_1_43
* net 89 wl_1_44
* net 90 wl_0_44
* net 91 wl_0_45
* net 92 wl_1_45
* net 93 wl_1_46
* net 94 wl_0_46
* net 95 wl_0_47
* net 96 wl_1_47
* net 97 wl_1_48
* net 98 wl_0_48
* net 99 wl_0_49
* net 100 wl_1_49
* net 101 wl_1_50
* net 102 wl_0_50
* net 103 wl_0_51
* net 104 wl_1_51
* net 105 wl_1_52
* net 106 wl_0_52
* net 107 wl_0_53
* net 108 wl_1_53
* net 109 wl_1_54
* net 110 wl_0_54
* net 111 wl_0_55
* net 112 wl_1_55
* net 113 wl_1_56
* net 114 wl_0_56
* net 115 wl_0_57
* net 116 wl_1_57
* net 117 wl_1_58
* net 118 wl_0_58
* net 119 wl_0_59
* net 120 wl_1_59
* net 121 wl_1_60
* net 122 wl_0_60
* net 123 wl_0_61
* net 124 wl_1_61
* net 125 wl_1_62
* net 126 wl_0_62
* net 127 wl_0_63
* net 128 wl_1_63
* net 129 wl_1_64
* net 130 wl_0_64
* net 131 wl_0_65
* net 132 wl_1_65
* net 133 wl_1_66
* net 134 wl_0_66
* net 135 wl_0_67
* net 136 wl_1_67
* net 137 vdd
* net 138 gnd
* cell instance $1 r0 *1 0,0
X$1 1 2 137 138 dummy_cell_2rw
* cell instance $2 m0 *1 0,2.99
X$2 4 3 137 138 dummy_cell_2rw
* cell instance $3 r0 *1 0,2.99
X$3 5 6 137 138 dummy_cell_2rw
* cell instance $4 m0 *1 0,5.98
X$4 8 7 137 138 dummy_cell_2rw
* cell instance $5 r0 *1 0,5.98
X$5 9 10 137 138 dummy_cell_2rw
* cell instance $6 m0 *1 0,8.97
X$6 12 11 137 138 dummy_cell_2rw
* cell instance $7 r0 *1 0,8.97
X$7 13 14 137 138 dummy_cell_2rw
* cell instance $8 m0 *1 0,11.96
X$8 16 15 137 138 dummy_cell_2rw
* cell instance $9 r0 *1 0,11.96
X$9 17 18 137 138 dummy_cell_2rw
* cell instance $10 m0 *1 0,14.95
X$10 20 19 137 138 dummy_cell_2rw
* cell instance $11 r0 *1 0,14.95
X$11 21 22 137 138 dummy_cell_2rw
* cell instance $12 m0 *1 0,17.94
X$12 24 23 137 138 dummy_cell_2rw
* cell instance $13 r0 *1 0,17.94
X$13 25 26 137 138 dummy_cell_2rw
* cell instance $14 m0 *1 0,20.93
X$14 28 27 137 138 dummy_cell_2rw
* cell instance $15 r0 *1 0,20.93
X$15 29 30 137 138 dummy_cell_2rw
* cell instance $16 m0 *1 0,23.92
X$16 32 31 137 138 dummy_cell_2rw
* cell instance $17 r0 *1 0,23.92
X$17 33 34 137 138 dummy_cell_2rw
* cell instance $18 m0 *1 0,26.91
X$18 36 35 137 138 dummy_cell_2rw
* cell instance $19 r0 *1 0,26.91
X$19 37 38 137 138 dummy_cell_2rw
* cell instance $20 m0 *1 0,29.9
X$20 40 39 137 138 dummy_cell_2rw
* cell instance $21 r0 *1 0,29.9
X$21 41 42 137 138 dummy_cell_2rw
* cell instance $22 m0 *1 0,32.89
X$22 44 43 137 138 dummy_cell_2rw
* cell instance $23 r0 *1 0,32.89
X$23 45 46 137 138 dummy_cell_2rw
* cell instance $24 m0 *1 0,35.88
X$24 48 47 137 138 dummy_cell_2rw
* cell instance $25 r0 *1 0,35.88
X$25 49 50 137 138 dummy_cell_2rw
* cell instance $26 m0 *1 0,38.87
X$26 52 51 137 138 dummy_cell_2rw
* cell instance $27 r0 *1 0,38.87
X$27 53 54 137 138 dummy_cell_2rw
* cell instance $28 m0 *1 0,41.86
X$28 56 55 137 138 dummy_cell_2rw
* cell instance $29 r0 *1 0,41.86
X$29 57 58 137 138 dummy_cell_2rw
* cell instance $30 m0 *1 0,44.85
X$30 60 59 137 138 dummy_cell_2rw
* cell instance $31 r0 *1 0,44.85
X$31 61 62 137 138 dummy_cell_2rw
* cell instance $32 m0 *1 0,47.84
X$32 64 63 137 138 dummy_cell_2rw
* cell instance $33 r0 *1 0,47.84
X$33 65 66 137 138 dummy_cell_2rw
* cell instance $34 m0 *1 0,50.83
X$34 68 67 137 138 dummy_cell_2rw
* cell instance $35 r0 *1 0,50.83
X$35 69 70 137 138 dummy_cell_2rw
* cell instance $36 m0 *1 0,53.82
X$36 72 71 137 138 dummy_cell_2rw
* cell instance $37 r0 *1 0,53.82
X$37 73 74 137 138 dummy_cell_2rw
* cell instance $38 m0 *1 0,56.81
X$38 76 75 137 138 dummy_cell_2rw
* cell instance $39 r0 *1 0,56.81
X$39 77 78 137 138 dummy_cell_2rw
* cell instance $40 m0 *1 0,59.8
X$40 80 79 137 138 dummy_cell_2rw
* cell instance $41 r0 *1 0,59.8
X$41 81 82 137 138 dummy_cell_2rw
* cell instance $42 m0 *1 0,62.79
X$42 84 83 137 138 dummy_cell_2rw
* cell instance $43 r0 *1 0,62.79
X$43 85 86 137 138 dummy_cell_2rw
* cell instance $44 m0 *1 0,65.78
X$44 88 87 137 138 dummy_cell_2rw
* cell instance $45 r0 *1 0,65.78
X$45 89 90 137 138 dummy_cell_2rw
* cell instance $46 m0 *1 0,68.77
X$46 92 91 137 138 dummy_cell_2rw
* cell instance $47 r0 *1 0,68.77
X$47 93 94 137 138 dummy_cell_2rw
* cell instance $48 m0 *1 0,71.76
X$48 96 95 137 138 dummy_cell_2rw
* cell instance $49 r0 *1 0,71.76
X$49 97 98 137 138 dummy_cell_2rw
* cell instance $50 m0 *1 0,74.75
X$50 100 99 137 138 dummy_cell_2rw
* cell instance $51 r0 *1 0,74.75
X$51 101 102 137 138 dummy_cell_2rw
* cell instance $52 m0 *1 0,77.74
X$52 104 103 137 138 dummy_cell_2rw
* cell instance $53 r0 *1 0,77.74
X$53 105 106 137 138 dummy_cell_2rw
* cell instance $54 m0 *1 0,80.73
X$54 108 107 137 138 dummy_cell_2rw
* cell instance $55 r0 *1 0,80.73
X$55 109 110 137 138 dummy_cell_2rw
* cell instance $56 m0 *1 0,83.72
X$56 112 111 137 138 dummy_cell_2rw
* cell instance $57 r0 *1 0,83.72
X$57 113 114 137 138 dummy_cell_2rw
* cell instance $58 m0 *1 0,86.71
X$58 116 115 137 138 dummy_cell_2rw
* cell instance $59 r0 *1 0,86.71
X$59 117 118 137 138 dummy_cell_2rw
* cell instance $60 m0 *1 0,89.7
X$60 120 119 137 138 dummy_cell_2rw
* cell instance $61 r0 *1 0,89.7
X$61 121 122 137 138 dummy_cell_2rw
* cell instance $62 m0 *1 0,92.69
X$62 124 123 137 138 dummy_cell_2rw
* cell instance $63 r0 *1 0,92.69
X$63 125 126 137 138 dummy_cell_2rw
* cell instance $64 m0 *1 0,95.68
X$64 128 127 137 138 dummy_cell_2rw
* cell instance $65 r0 *1 0,95.68
X$65 129 130 137 138 dummy_cell_2rw
* cell instance $66 m0 *1 0,98.67
X$66 132 131 137 138 dummy_cell_2rw
* cell instance $67 r0 *1 0,98.67
X$67 133 134 137 138 dummy_cell_2rw
* cell instance $68 m0 *1 0,101.66
X$68 136 135 137 138 dummy_cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_dummy_array_3

* cell custom_sram_1r1w_32_256_freepdk45_dummy_array_2
* pin wl_1_0
* pin wl_0_0
* pin wl_0_1
* pin wl_1_1
* pin wl_1_2
* pin wl_0_2
* pin wl_0_3
* pin wl_1_3
* pin wl_1_4
* pin wl_0_4
* pin wl_0_5
* pin wl_1_5
* pin wl_1_6
* pin wl_0_6
* pin wl_0_7
* pin wl_1_7
* pin wl_1_8
* pin wl_0_8
* pin wl_0_9
* pin wl_1_9
* pin wl_1_10
* pin wl_0_10
* pin wl_0_11
* pin wl_1_11
* pin wl_1_12
* pin wl_0_12
* pin wl_0_13
* pin wl_1_13
* pin wl_1_14
* pin wl_0_14
* pin wl_0_15
* pin wl_1_15
* pin wl_1_16
* pin wl_0_16
* pin wl_0_17
* pin wl_1_17
* pin wl_1_18
* pin wl_0_18
* pin wl_0_19
* pin wl_1_19
* pin wl_1_20
* pin wl_0_20
* pin wl_0_21
* pin wl_1_21
* pin wl_1_22
* pin wl_0_22
* pin wl_0_23
* pin wl_1_23
* pin wl_1_24
* pin wl_0_24
* pin wl_0_25
* pin wl_1_25
* pin wl_1_26
* pin wl_0_26
* pin wl_0_27
* pin wl_1_27
* pin wl_1_28
* pin wl_0_28
* pin wl_0_29
* pin wl_1_29
* pin wl_1_30
* pin wl_0_30
* pin wl_0_31
* pin wl_1_31
* pin wl_1_32
* pin wl_0_32
* pin wl_0_33
* pin wl_1_33
* pin wl_1_34
* pin wl_0_34
* pin wl_0_35
* pin wl_1_35
* pin wl_1_36
* pin wl_0_36
* pin wl_0_37
* pin wl_1_37
* pin wl_1_38
* pin wl_0_38
* pin wl_0_39
* pin wl_1_39
* pin wl_1_40
* pin wl_0_40
* pin wl_0_41
* pin wl_1_41
* pin wl_1_42
* pin wl_0_42
* pin wl_0_43
* pin wl_1_43
* pin wl_1_44
* pin wl_0_44
* pin wl_0_45
* pin wl_1_45
* pin wl_1_46
* pin wl_0_46
* pin wl_0_47
* pin wl_1_47
* pin wl_1_48
* pin wl_0_48
* pin wl_0_49
* pin wl_1_49
* pin wl_1_50
* pin wl_0_50
* pin wl_0_51
* pin wl_1_51
* pin wl_1_52
* pin wl_0_52
* pin wl_0_53
* pin wl_1_53
* pin wl_1_54
* pin wl_0_54
* pin wl_0_55
* pin wl_1_55
* pin wl_1_56
* pin wl_0_56
* pin wl_0_57
* pin wl_1_57
* pin wl_1_58
* pin wl_0_58
* pin wl_0_59
* pin wl_1_59
* pin wl_1_60
* pin wl_0_60
* pin wl_0_61
* pin wl_1_61
* pin wl_1_62
* pin wl_0_62
* pin wl_0_63
* pin wl_1_63
* pin wl_1_64
* pin wl_0_64
* pin wl_0_65
* pin wl_1_65
* pin wl_1_66
* pin wl_0_66
* pin wl_0_67
* pin wl_1_67
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_dummy_array_2 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37
+ 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89
+ 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111
+ 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130
+ 131 132 133 134 135 136 137 138
* net 1 wl_1_0
* net 2 wl_0_0
* net 3 wl_0_1
* net 4 wl_1_1
* net 5 wl_1_2
* net 6 wl_0_2
* net 7 wl_0_3
* net 8 wl_1_3
* net 9 wl_1_4
* net 10 wl_0_4
* net 11 wl_0_5
* net 12 wl_1_5
* net 13 wl_1_6
* net 14 wl_0_6
* net 15 wl_0_7
* net 16 wl_1_7
* net 17 wl_1_8
* net 18 wl_0_8
* net 19 wl_0_9
* net 20 wl_1_9
* net 21 wl_1_10
* net 22 wl_0_10
* net 23 wl_0_11
* net 24 wl_1_11
* net 25 wl_1_12
* net 26 wl_0_12
* net 27 wl_0_13
* net 28 wl_1_13
* net 29 wl_1_14
* net 30 wl_0_14
* net 31 wl_0_15
* net 32 wl_1_15
* net 33 wl_1_16
* net 34 wl_0_16
* net 35 wl_0_17
* net 36 wl_1_17
* net 37 wl_1_18
* net 38 wl_0_18
* net 39 wl_0_19
* net 40 wl_1_19
* net 41 wl_1_20
* net 42 wl_0_20
* net 43 wl_0_21
* net 44 wl_1_21
* net 45 wl_1_22
* net 46 wl_0_22
* net 47 wl_0_23
* net 48 wl_1_23
* net 49 wl_1_24
* net 50 wl_0_24
* net 51 wl_0_25
* net 52 wl_1_25
* net 53 wl_1_26
* net 54 wl_0_26
* net 55 wl_0_27
* net 56 wl_1_27
* net 57 wl_1_28
* net 58 wl_0_28
* net 59 wl_0_29
* net 60 wl_1_29
* net 61 wl_1_30
* net 62 wl_0_30
* net 63 wl_0_31
* net 64 wl_1_31
* net 65 wl_1_32
* net 66 wl_0_32
* net 67 wl_0_33
* net 68 wl_1_33
* net 69 wl_1_34
* net 70 wl_0_34
* net 71 wl_0_35
* net 72 wl_1_35
* net 73 wl_1_36
* net 74 wl_0_36
* net 75 wl_0_37
* net 76 wl_1_37
* net 77 wl_1_38
* net 78 wl_0_38
* net 79 wl_0_39
* net 80 wl_1_39
* net 81 wl_1_40
* net 82 wl_0_40
* net 83 wl_0_41
* net 84 wl_1_41
* net 85 wl_1_42
* net 86 wl_0_42
* net 87 wl_0_43
* net 88 wl_1_43
* net 89 wl_1_44
* net 90 wl_0_44
* net 91 wl_0_45
* net 92 wl_1_45
* net 93 wl_1_46
* net 94 wl_0_46
* net 95 wl_0_47
* net 96 wl_1_47
* net 97 wl_1_48
* net 98 wl_0_48
* net 99 wl_0_49
* net 100 wl_1_49
* net 101 wl_1_50
* net 102 wl_0_50
* net 103 wl_0_51
* net 104 wl_1_51
* net 105 wl_1_52
* net 106 wl_0_52
* net 107 wl_0_53
* net 108 wl_1_53
* net 109 wl_1_54
* net 110 wl_0_54
* net 111 wl_0_55
* net 112 wl_1_55
* net 113 wl_1_56
* net 114 wl_0_56
* net 115 wl_0_57
* net 116 wl_1_57
* net 117 wl_1_58
* net 118 wl_0_58
* net 119 wl_0_59
* net 120 wl_1_59
* net 121 wl_1_60
* net 122 wl_0_60
* net 123 wl_0_61
* net 124 wl_1_61
* net 125 wl_1_62
* net 126 wl_0_62
* net 127 wl_0_63
* net 128 wl_1_63
* net 129 wl_1_64
* net 130 wl_0_64
* net 131 wl_0_65
* net 132 wl_1_65
* net 133 wl_1_66
* net 134 wl_0_66
* net 135 wl_0_67
* net 136 wl_1_67
* net 137 vdd
* net 138 gnd
* cell instance $1 r0 *1 0,0
X$1 1 2 137 138 dummy_cell_2rw
* cell instance $2 m0 *1 0,2.99
X$2 4 3 137 138 dummy_cell_2rw
* cell instance $3 r0 *1 0,2.99
X$3 5 6 137 138 dummy_cell_2rw
* cell instance $4 m0 *1 0,5.98
X$4 8 7 137 138 dummy_cell_2rw
* cell instance $5 r0 *1 0,5.98
X$5 9 10 137 138 dummy_cell_2rw
* cell instance $6 m0 *1 0,8.97
X$6 12 11 137 138 dummy_cell_2rw
* cell instance $7 r0 *1 0,8.97
X$7 13 14 137 138 dummy_cell_2rw
* cell instance $8 m0 *1 0,11.96
X$8 16 15 137 138 dummy_cell_2rw
* cell instance $9 r0 *1 0,11.96
X$9 17 18 137 138 dummy_cell_2rw
* cell instance $10 m0 *1 0,14.95
X$10 20 19 137 138 dummy_cell_2rw
* cell instance $11 r0 *1 0,14.95
X$11 21 22 137 138 dummy_cell_2rw
* cell instance $12 m0 *1 0,17.94
X$12 24 23 137 138 dummy_cell_2rw
* cell instance $13 r0 *1 0,17.94
X$13 25 26 137 138 dummy_cell_2rw
* cell instance $14 m0 *1 0,20.93
X$14 28 27 137 138 dummy_cell_2rw
* cell instance $15 r0 *1 0,20.93
X$15 29 30 137 138 dummy_cell_2rw
* cell instance $16 m0 *1 0,23.92
X$16 32 31 137 138 dummy_cell_2rw
* cell instance $17 r0 *1 0,23.92
X$17 33 34 137 138 dummy_cell_2rw
* cell instance $18 m0 *1 0,26.91
X$18 36 35 137 138 dummy_cell_2rw
* cell instance $19 r0 *1 0,26.91
X$19 37 38 137 138 dummy_cell_2rw
* cell instance $20 m0 *1 0,29.9
X$20 40 39 137 138 dummy_cell_2rw
* cell instance $21 r0 *1 0,29.9
X$21 41 42 137 138 dummy_cell_2rw
* cell instance $22 m0 *1 0,32.89
X$22 44 43 137 138 dummy_cell_2rw
* cell instance $23 r0 *1 0,32.89
X$23 45 46 137 138 dummy_cell_2rw
* cell instance $24 m0 *1 0,35.88
X$24 48 47 137 138 dummy_cell_2rw
* cell instance $25 r0 *1 0,35.88
X$25 49 50 137 138 dummy_cell_2rw
* cell instance $26 m0 *1 0,38.87
X$26 52 51 137 138 dummy_cell_2rw
* cell instance $27 r0 *1 0,38.87
X$27 53 54 137 138 dummy_cell_2rw
* cell instance $28 m0 *1 0,41.86
X$28 56 55 137 138 dummy_cell_2rw
* cell instance $29 r0 *1 0,41.86
X$29 57 58 137 138 dummy_cell_2rw
* cell instance $30 m0 *1 0,44.85
X$30 60 59 137 138 dummy_cell_2rw
* cell instance $31 r0 *1 0,44.85
X$31 61 62 137 138 dummy_cell_2rw
* cell instance $32 m0 *1 0,47.84
X$32 64 63 137 138 dummy_cell_2rw
* cell instance $33 r0 *1 0,47.84
X$33 65 66 137 138 dummy_cell_2rw
* cell instance $34 m0 *1 0,50.83
X$34 68 67 137 138 dummy_cell_2rw
* cell instance $35 r0 *1 0,50.83
X$35 69 70 137 138 dummy_cell_2rw
* cell instance $36 m0 *1 0,53.82
X$36 72 71 137 138 dummy_cell_2rw
* cell instance $37 r0 *1 0,53.82
X$37 73 74 137 138 dummy_cell_2rw
* cell instance $38 m0 *1 0,56.81
X$38 76 75 137 138 dummy_cell_2rw
* cell instance $39 r0 *1 0,56.81
X$39 77 78 137 138 dummy_cell_2rw
* cell instance $40 m0 *1 0,59.8
X$40 80 79 137 138 dummy_cell_2rw
* cell instance $41 r0 *1 0,59.8
X$41 81 82 137 138 dummy_cell_2rw
* cell instance $42 m0 *1 0,62.79
X$42 84 83 137 138 dummy_cell_2rw
* cell instance $43 r0 *1 0,62.79
X$43 85 86 137 138 dummy_cell_2rw
* cell instance $44 m0 *1 0,65.78
X$44 88 87 137 138 dummy_cell_2rw
* cell instance $45 r0 *1 0,65.78
X$45 89 90 137 138 dummy_cell_2rw
* cell instance $46 m0 *1 0,68.77
X$46 92 91 137 138 dummy_cell_2rw
* cell instance $47 r0 *1 0,68.77
X$47 93 94 137 138 dummy_cell_2rw
* cell instance $48 m0 *1 0,71.76
X$48 96 95 137 138 dummy_cell_2rw
* cell instance $49 r0 *1 0,71.76
X$49 97 98 137 138 dummy_cell_2rw
* cell instance $50 m0 *1 0,74.75
X$50 100 99 137 138 dummy_cell_2rw
* cell instance $51 r0 *1 0,74.75
X$51 101 102 137 138 dummy_cell_2rw
* cell instance $52 m0 *1 0,77.74
X$52 104 103 137 138 dummy_cell_2rw
* cell instance $53 r0 *1 0,77.74
X$53 105 106 137 138 dummy_cell_2rw
* cell instance $54 m0 *1 0,80.73
X$54 108 107 137 138 dummy_cell_2rw
* cell instance $55 r0 *1 0,80.73
X$55 109 110 137 138 dummy_cell_2rw
* cell instance $56 m0 *1 0,83.72
X$56 112 111 137 138 dummy_cell_2rw
* cell instance $57 r0 *1 0,83.72
X$57 113 114 137 138 dummy_cell_2rw
* cell instance $58 m0 *1 0,86.71
X$58 116 115 137 138 dummy_cell_2rw
* cell instance $59 r0 *1 0,86.71
X$59 117 118 137 138 dummy_cell_2rw
* cell instance $60 m0 *1 0,89.7
X$60 120 119 137 138 dummy_cell_2rw
* cell instance $61 r0 *1 0,89.7
X$61 121 122 137 138 dummy_cell_2rw
* cell instance $62 m0 *1 0,92.69
X$62 124 123 137 138 dummy_cell_2rw
* cell instance $63 r0 *1 0,92.69
X$63 125 126 137 138 dummy_cell_2rw
* cell instance $64 m0 *1 0,95.68
X$64 128 127 137 138 dummy_cell_2rw
* cell instance $65 r0 *1 0,95.68
X$65 129 130 137 138 dummy_cell_2rw
* cell instance $66 m0 *1 0,98.67
X$66 132 131 137 138 dummy_cell_2rw
* cell instance $67 r0 *1 0,98.67
X$67 133 134 137 138 dummy_cell_2rw
* cell instance $68 m0 *1 0,101.66
X$68 136 135 137 138 dummy_cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_dummy_array_2

* cell custom_sram_1r1w_32_256_freepdk45_dummy_array_0
* pin wl_0_0
* pin wl_1_0
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_dummy_array_0 1 2 3 4
* net 1 wl_0_0
* net 2 wl_1_0
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 dummy_cell_2rw
* cell instance $2 r0 *1 1.175,0
X$2 2 1 3 4 dummy_cell_2rw
* cell instance $3 r0 *1 2.35,0
X$3 2 1 3 4 dummy_cell_2rw
* cell instance $4 r0 *1 3.525,0
X$4 2 1 3 4 dummy_cell_2rw
* cell instance $5 r0 *1 4.7,0
X$5 2 1 3 4 dummy_cell_2rw
* cell instance $6 r0 *1 5.875,0
X$6 2 1 3 4 dummy_cell_2rw
* cell instance $7 r0 *1 7.05,0
X$7 2 1 3 4 dummy_cell_2rw
* cell instance $8 r0 *1 8.225,0
X$8 2 1 3 4 dummy_cell_2rw
* cell instance $9 r0 *1 9.4,0
X$9 2 1 3 4 dummy_cell_2rw
* cell instance $10 r0 *1 10.575,0
X$10 2 1 3 4 dummy_cell_2rw
* cell instance $11 r0 *1 11.75,0
X$11 2 1 3 4 dummy_cell_2rw
* cell instance $12 r0 *1 12.925,0
X$12 2 1 3 4 dummy_cell_2rw
* cell instance $13 r0 *1 14.1,0
X$13 2 1 3 4 dummy_cell_2rw
* cell instance $14 r0 *1 15.275,0
X$14 2 1 3 4 dummy_cell_2rw
* cell instance $15 r0 *1 16.45,0
X$15 2 1 3 4 dummy_cell_2rw
* cell instance $16 r0 *1 17.625,0
X$16 2 1 3 4 dummy_cell_2rw
* cell instance $17 r0 *1 18.8,0
X$17 2 1 3 4 dummy_cell_2rw
* cell instance $18 r0 *1 19.975,0
X$18 2 1 3 4 dummy_cell_2rw
* cell instance $19 r0 *1 21.15,0
X$19 2 1 3 4 dummy_cell_2rw
* cell instance $20 r0 *1 22.325,0
X$20 2 1 3 4 dummy_cell_2rw
* cell instance $21 r0 *1 23.5,0
X$21 2 1 3 4 dummy_cell_2rw
* cell instance $22 r0 *1 24.675,0
X$22 2 1 3 4 dummy_cell_2rw
* cell instance $23 r0 *1 25.85,0
X$23 2 1 3 4 dummy_cell_2rw
* cell instance $24 r0 *1 27.025,0
X$24 2 1 3 4 dummy_cell_2rw
* cell instance $25 r0 *1 28.2,0
X$25 2 1 3 4 dummy_cell_2rw
* cell instance $26 r0 *1 29.375,0
X$26 2 1 3 4 dummy_cell_2rw
* cell instance $27 r0 *1 30.55,0
X$27 2 1 3 4 dummy_cell_2rw
* cell instance $28 r0 *1 31.725,0
X$28 2 1 3 4 dummy_cell_2rw
* cell instance $29 r0 *1 32.9,0
X$29 2 1 3 4 dummy_cell_2rw
* cell instance $30 r0 *1 34.075,0
X$30 2 1 3 4 dummy_cell_2rw
* cell instance $31 r0 *1 35.25,0
X$31 2 1 3 4 dummy_cell_2rw
* cell instance $32 r0 *1 36.425,0
X$32 2 1 3 4 dummy_cell_2rw
* cell instance $33 r0 *1 37.6,0
X$33 2 1 3 4 dummy_cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_dummy_array_0

* cell custom_sram_1r1w_32_256_freepdk45_dummy_array_1
* pin wl_0_0
* pin wl_1_0
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_dummy_array_1 1 2 3 4
* net 1 wl_0_0
* net 2 wl_1_0
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 dummy_cell_2rw
* cell instance $2 r0 *1 1.175,0
X$2 2 1 3 4 dummy_cell_2rw
* cell instance $3 r0 *1 2.35,0
X$3 2 1 3 4 dummy_cell_2rw
* cell instance $4 r0 *1 3.525,0
X$4 2 1 3 4 dummy_cell_2rw
* cell instance $5 r0 *1 4.7,0
X$5 2 1 3 4 dummy_cell_2rw
* cell instance $6 r0 *1 5.875,0
X$6 2 1 3 4 dummy_cell_2rw
* cell instance $7 r0 *1 7.05,0
X$7 2 1 3 4 dummy_cell_2rw
* cell instance $8 r0 *1 8.225,0
X$8 2 1 3 4 dummy_cell_2rw
* cell instance $9 r0 *1 9.4,0
X$9 2 1 3 4 dummy_cell_2rw
* cell instance $10 r0 *1 10.575,0
X$10 2 1 3 4 dummy_cell_2rw
* cell instance $11 r0 *1 11.75,0
X$11 2 1 3 4 dummy_cell_2rw
* cell instance $12 r0 *1 12.925,0
X$12 2 1 3 4 dummy_cell_2rw
* cell instance $13 r0 *1 14.1,0
X$13 2 1 3 4 dummy_cell_2rw
* cell instance $14 r0 *1 15.275,0
X$14 2 1 3 4 dummy_cell_2rw
* cell instance $15 r0 *1 16.45,0
X$15 2 1 3 4 dummy_cell_2rw
* cell instance $16 r0 *1 17.625,0
X$16 2 1 3 4 dummy_cell_2rw
* cell instance $17 r0 *1 18.8,0
X$17 2 1 3 4 dummy_cell_2rw
* cell instance $18 r0 *1 19.975,0
X$18 2 1 3 4 dummy_cell_2rw
* cell instance $19 r0 *1 21.15,0
X$19 2 1 3 4 dummy_cell_2rw
* cell instance $20 r0 *1 22.325,0
X$20 2 1 3 4 dummy_cell_2rw
* cell instance $21 r0 *1 23.5,0
X$21 2 1 3 4 dummy_cell_2rw
* cell instance $22 r0 *1 24.675,0
X$22 2 1 3 4 dummy_cell_2rw
* cell instance $23 r0 *1 25.85,0
X$23 2 1 3 4 dummy_cell_2rw
* cell instance $24 r0 *1 27.025,0
X$24 2 1 3 4 dummy_cell_2rw
* cell instance $25 r0 *1 28.2,0
X$25 2 1 3 4 dummy_cell_2rw
* cell instance $26 r0 *1 29.375,0
X$26 2 1 3 4 dummy_cell_2rw
* cell instance $27 r0 *1 30.55,0
X$27 2 1 3 4 dummy_cell_2rw
* cell instance $28 r0 *1 31.725,0
X$28 2 1 3 4 dummy_cell_2rw
* cell instance $29 r0 *1 32.9,0
X$29 2 1 3 4 dummy_cell_2rw
* cell instance $30 r0 *1 34.075,0
X$30 2 1 3 4 dummy_cell_2rw
* cell instance $31 r0 *1 35.25,0
X$31 2 1 3 4 dummy_cell_2rw
* cell instance $32 r0 *1 36.425,0
X$32 2 1 3 4 dummy_cell_2rw
* cell instance $33 r0 *1 37.6,0
X$33 2 1 3 4 dummy_cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_dummy_array_1

* cell custom_sram_1r1w_32_256_freepdk45_replica_bitcell_array
* pin rbl_wl_0_0
* pin rbl_wl_0_1
* pin rbl_bl_0_0
* pin rbl_bl_1_0
* pin rbl_br_1_0
* pin rbl_br_0_0
* pin bl_0_0
* pin bl_1_0
* pin br_1_0
* pin br_0_0
* pin bl_0_1
* pin bl_1_1
* pin br_1_1
* pin br_0_1
* pin bl_0_2
* pin bl_1_2
* pin br_1_2
* pin br_0_2
* pin bl_0_3
* pin bl_1_3
* pin br_1_3
* pin br_0_3
* pin bl_0_4
* pin bl_1_4
* pin br_1_4
* pin br_0_4
* pin bl_0_5
* pin bl_1_5
* pin br_1_5
* pin br_0_5
* pin bl_0_6
* pin bl_1_6
* pin br_1_6
* pin br_0_6
* pin bl_0_7
* pin bl_1_7
* pin br_1_7
* pin br_0_7
* pin bl_0_8
* pin bl_1_8
* pin br_1_8
* pin br_0_8
* pin bl_0_9
* pin bl_1_9
* pin br_1_9
* pin br_0_9
* pin bl_0_10
* pin bl_1_10
* pin br_1_10
* pin br_0_10
* pin bl_0_11
* pin bl_1_11
* pin br_1_11
* pin br_0_11
* pin bl_0_12
* pin bl_1_12
* pin br_1_12
* pin br_0_12
* pin bl_0_13
* pin bl_1_13
* pin br_1_13
* pin br_0_13
* pin bl_0_14
* pin bl_1_14
* pin br_1_14
* pin br_0_14
* pin bl_0_15
* pin bl_1_15
* pin br_1_15
* pin br_0_15
* pin bl_0_16
* pin bl_1_16
* pin br_1_16
* pin br_0_16
* pin bl_0_17
* pin bl_1_17
* pin br_1_17
* pin br_0_17
* pin bl_0_18
* pin bl_1_18
* pin br_1_18
* pin br_0_18
* pin bl_0_19
* pin bl_1_19
* pin br_1_19
* pin br_0_19
* pin bl_0_20
* pin bl_1_20
* pin br_1_20
* pin br_0_20
* pin bl_0_21
* pin bl_1_21
* pin br_1_21
* pin br_0_21
* pin bl_0_22
* pin bl_1_22
* pin br_1_22
* pin br_0_22
* pin bl_0_23
* pin bl_1_23
* pin br_1_23
* pin br_0_23
* pin bl_0_24
* pin bl_1_24
* pin br_1_24
* pin br_0_24
* pin bl_0_25
* pin bl_1_25
* pin br_1_25
* pin br_0_25
* pin bl_0_26
* pin bl_1_26
* pin br_1_26
* pin br_0_26
* pin bl_0_27
* pin bl_1_27
* pin br_1_27
* pin br_0_27
* pin bl_0_28
* pin bl_1_28
* pin br_1_28
* pin br_0_28
* pin bl_0_29
* pin bl_1_29
* pin br_1_29
* pin br_0_29
* pin bl_0_30
* pin bl_1_30
* pin br_1_30
* pin br_0_30
* pin bl_0_31
* pin bl_1_31
* pin br_1_31
* pin br_0_31
* pin wl_1_0
* pin wl_0_0
* pin wl_1_1
* pin wl_0_1
* pin wl_0_2
* pin wl_1_2
* pin wl_1_3
* pin wl_0_3
* pin wl_0_4
* pin wl_1_4
* pin wl_1_5
* pin wl_0_5
* pin wl_0_6
* pin wl_1_6
* pin wl_0_7
* pin wl_1_7
* pin wl_0_8
* pin wl_1_8
* pin wl_0_9
* pin wl_1_9
* pin wl_0_10
* pin wl_1_10
* pin wl_1_11
* pin wl_0_11
* pin wl_0_12
* pin wl_1_12
* pin wl_1_13
* pin wl_0_13
* pin wl_0_14
* pin wl_1_14
* pin wl_1_15
* pin wl_0_15
* pin wl_0_16
* pin wl_1_16
* pin wl_1_17
* pin wl_0_17
* pin wl_0_18
* pin wl_1_18
* pin wl_1_19
* pin wl_0_19
* pin wl_0_20
* pin wl_1_20
* pin wl_1_21
* pin wl_0_21
* pin wl_1_22
* pin wl_0_22
* pin wl_0_23
* pin wl_1_23
* pin wl_1_24
* pin wl_0_24
* pin wl_1_25
* pin wl_0_25
* pin wl_0_26
* pin wl_1_26
* pin wl_1_27
* pin wl_0_27
* pin wl_0_28
* pin wl_1_28
* pin wl_1_29
* pin wl_0_29
* pin wl_0_30
* pin wl_1_30
* pin wl_1_31
* pin wl_0_31
* pin wl_1_32
* pin wl_0_32
* pin wl_1_33
* pin wl_0_33
* pin wl_0_34
* pin wl_1_34
* pin wl_1_35
* pin wl_0_35
* pin wl_0_36
* pin wl_1_36
* pin wl_0_37
* pin wl_1_37
* pin wl_0_38
* pin wl_1_38
* pin wl_0_39
* pin wl_1_39
* pin wl_0_40
* pin wl_1_40
* pin wl_1_41
* pin wl_0_41
* pin wl_0_42
* pin wl_1_42
* pin wl_1_43
* pin wl_0_43
* pin wl_0_44
* pin wl_1_44
* pin wl_1_45
* pin wl_0_45
* pin wl_0_46
* pin wl_1_46
* pin wl_1_47
* pin wl_0_47
* pin wl_0_48
* pin wl_1_48
* pin wl_0_49
* pin wl_1_49
* pin wl_0_50
* pin wl_1_50
* pin wl_1_51
* pin wl_0_51
* pin wl_0_52
* pin wl_1_52
* pin wl_1_53
* pin wl_0_53
* pin wl_1_54
* pin wl_0_54
* pin wl_1_55
* pin wl_0_55
* pin wl_1_56
* pin wl_0_56
* pin wl_1_57
* pin wl_0_57
* pin wl_1_58
* pin wl_0_58
* pin wl_1_59
* pin wl_0_59
* pin wl_0_60
* pin wl_1_60
* pin wl_0_61
* pin wl_1_61
* pin wl_1_62
* pin wl_0_62
* pin wl_0_63
* pin wl_1_63
* pin rbl_wl_1_1
* pin rbl_wl_1_0
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_replica_bitcell_array 1 2 3 4 5 6 7 8
+ 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34
+ 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86
+ 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108
+ 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127
+ 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146
+ 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165
+ 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184
+ 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266
* net 1 rbl_wl_0_0
* net 2 rbl_wl_0_1
* net 3 rbl_bl_0_0
* net 4 rbl_bl_1_0
* net 5 rbl_br_1_0
* net 6 rbl_br_0_0
* net 7 bl_0_0
* net 8 bl_1_0
* net 9 br_1_0
* net 10 br_0_0
* net 11 bl_0_1
* net 12 bl_1_1
* net 13 br_1_1
* net 14 br_0_1
* net 15 bl_0_2
* net 16 bl_1_2
* net 17 br_1_2
* net 18 br_0_2
* net 19 bl_0_3
* net 20 bl_1_3
* net 21 br_1_3
* net 22 br_0_3
* net 23 bl_0_4
* net 24 bl_1_4
* net 25 br_1_4
* net 26 br_0_4
* net 27 bl_0_5
* net 28 bl_1_5
* net 29 br_1_5
* net 30 br_0_5
* net 31 bl_0_6
* net 32 bl_1_6
* net 33 br_1_6
* net 34 br_0_6
* net 35 bl_0_7
* net 36 bl_1_7
* net 37 br_1_7
* net 38 br_0_7
* net 39 bl_0_8
* net 40 bl_1_8
* net 41 br_1_8
* net 42 br_0_8
* net 43 bl_0_9
* net 44 bl_1_9
* net 45 br_1_9
* net 46 br_0_9
* net 47 bl_0_10
* net 48 bl_1_10
* net 49 br_1_10
* net 50 br_0_10
* net 51 bl_0_11
* net 52 bl_1_11
* net 53 br_1_11
* net 54 br_0_11
* net 55 bl_0_12
* net 56 bl_1_12
* net 57 br_1_12
* net 58 br_0_12
* net 59 bl_0_13
* net 60 bl_1_13
* net 61 br_1_13
* net 62 br_0_13
* net 63 bl_0_14
* net 64 bl_1_14
* net 65 br_1_14
* net 66 br_0_14
* net 67 bl_0_15
* net 68 bl_1_15
* net 69 br_1_15
* net 70 br_0_15
* net 71 bl_0_16
* net 72 bl_1_16
* net 73 br_1_16
* net 74 br_0_16
* net 75 bl_0_17
* net 76 bl_1_17
* net 77 br_1_17
* net 78 br_0_17
* net 79 bl_0_18
* net 80 bl_1_18
* net 81 br_1_18
* net 82 br_0_18
* net 83 bl_0_19
* net 84 bl_1_19
* net 85 br_1_19
* net 86 br_0_19
* net 87 bl_0_20
* net 88 bl_1_20
* net 89 br_1_20
* net 90 br_0_20
* net 91 bl_0_21
* net 92 bl_1_21
* net 93 br_1_21
* net 94 br_0_21
* net 95 bl_0_22
* net 96 bl_1_22
* net 97 br_1_22
* net 98 br_0_22
* net 99 bl_0_23
* net 100 bl_1_23
* net 101 br_1_23
* net 102 br_0_23
* net 103 bl_0_24
* net 104 bl_1_24
* net 105 br_1_24
* net 106 br_0_24
* net 107 bl_0_25
* net 108 bl_1_25
* net 109 br_1_25
* net 110 br_0_25
* net 111 bl_0_26
* net 112 bl_1_26
* net 113 br_1_26
* net 114 br_0_26
* net 115 bl_0_27
* net 116 bl_1_27
* net 117 br_1_27
* net 118 br_0_27
* net 119 bl_0_28
* net 120 bl_1_28
* net 121 br_1_28
* net 122 br_0_28
* net 123 bl_0_29
* net 124 bl_1_29
* net 125 br_1_29
* net 126 br_0_29
* net 127 bl_0_30
* net 128 bl_1_30
* net 129 br_1_30
* net 130 br_0_30
* net 131 bl_0_31
* net 132 bl_1_31
* net 133 br_1_31
* net 134 br_0_31
* net 135 wl_1_0
* net 136 wl_0_0
* net 137 wl_1_1
* net 138 wl_0_1
* net 139 wl_0_2
* net 140 wl_1_2
* net 141 wl_1_3
* net 142 wl_0_3
* net 143 wl_0_4
* net 144 wl_1_4
* net 145 wl_1_5
* net 146 wl_0_5
* net 147 wl_0_6
* net 148 wl_1_6
* net 149 wl_0_7
* net 150 wl_1_7
* net 151 wl_0_8
* net 152 wl_1_8
* net 153 wl_0_9
* net 154 wl_1_9
* net 155 wl_0_10
* net 156 wl_1_10
* net 157 wl_1_11
* net 158 wl_0_11
* net 159 wl_0_12
* net 160 wl_1_12
* net 161 wl_1_13
* net 162 wl_0_13
* net 163 wl_0_14
* net 164 wl_1_14
* net 165 wl_1_15
* net 166 wl_0_15
* net 167 wl_0_16
* net 168 wl_1_16
* net 169 wl_1_17
* net 170 wl_0_17
* net 171 wl_0_18
* net 172 wl_1_18
* net 173 wl_1_19
* net 174 wl_0_19
* net 175 wl_0_20
* net 176 wl_1_20
* net 177 wl_1_21
* net 178 wl_0_21
* net 179 wl_1_22
* net 180 wl_0_22
* net 181 wl_0_23
* net 182 wl_1_23
* net 183 wl_1_24
* net 184 wl_0_24
* net 185 wl_1_25
* net 186 wl_0_25
* net 187 wl_0_26
* net 188 wl_1_26
* net 189 wl_1_27
* net 190 wl_0_27
* net 191 wl_0_28
* net 192 wl_1_28
* net 193 wl_1_29
* net 194 wl_0_29
* net 195 wl_0_30
* net 196 wl_1_30
* net 197 wl_1_31
* net 198 wl_0_31
* net 199 wl_1_32
* net 200 wl_0_32
* net 201 wl_1_33
* net 202 wl_0_33
* net 203 wl_0_34
* net 204 wl_1_34
* net 205 wl_1_35
* net 206 wl_0_35
* net 207 wl_0_36
* net 208 wl_1_36
* net 209 wl_0_37
* net 210 wl_1_37
* net 211 wl_0_38
* net 212 wl_1_38
* net 213 wl_0_39
* net 214 wl_1_39
* net 215 wl_0_40
* net 216 wl_1_40
* net 217 wl_1_41
* net 218 wl_0_41
* net 219 wl_0_42
* net 220 wl_1_42
* net 221 wl_1_43
* net 222 wl_0_43
* net 223 wl_0_44
* net 224 wl_1_44
* net 225 wl_1_45
* net 226 wl_0_45
* net 227 wl_0_46
* net 228 wl_1_46
* net 229 wl_1_47
* net 230 wl_0_47
* net 231 wl_0_48
* net 232 wl_1_48
* net 233 wl_0_49
* net 234 wl_1_49
* net 235 wl_0_50
* net 236 wl_1_50
* net 237 wl_1_51
* net 238 wl_0_51
* net 239 wl_0_52
* net 240 wl_1_52
* net 241 wl_1_53
* net 242 wl_0_53
* net 243 wl_1_54
* net 244 wl_0_54
* net 245 wl_1_55
* net 246 wl_0_55
* net 247 wl_1_56
* net 248 wl_0_56
* net 249 wl_1_57
* net 250 wl_0_57
* net 251 wl_1_58
* net 252 wl_0_58
* net 253 wl_1_59
* net 254 wl_0_59
* net 255 wl_0_60
* net 256 wl_1_60
* net 257 wl_0_61
* net 258 wl_1_61
* net 259 wl_1_62
* net 260 wl_0_62
* net 261 wl_0_63
* net 262 wl_1_63
* net 263 rbl_wl_1_1
* net 264 rbl_wl_1_0
* net 265 vdd
* net 266 gnd
* cell instance $1 r0 *1 0,0
X$1 1 2 135 136 138 137 140 139 142 141 144 143 146 145 148 147 149 150 152 151
+ 153 154 156 155 158 157 160 159 162 161 164 163 166 165 168 167 170 169 172
+ 171 174 173 176 175 178 177 179 180 181 182 183 184 186 185 188 187 190 189
+ 192 191 194 193 196 195 3 4 198 197 5 6 199 200 202 201 204 203 206 205 208
+ 207 209 210 212 211 213 214 216 215 218 217 220 219 222 221 224 223 226 225
+ 228 227 230 229 232 231 233 234 236 235 238 237 240 239 242 241 243 244 246
+ 245 247 248 250 249 251 252 254 253 256 255 257 258 259 260 261 262 263 264
+ 265 266 custom_sram_1r1w_32_256_freepdk45_replica_column
* cell instance $2 m0 *1 1.175,1.495
X$2 1 2 265 266 custom_sram_1r1w_32_256_freepdk45_dummy_array
* cell instance $3 r0 *1 1.175,1.495
X$3 139 140 138 137 136 135 144 146 145 143 141 142 150 149 151 152 148 147 155
+ 156 157 158 153 154 163 161 160 164 162 159 168 170 167 169 165 166 176 175
+ 171 174 173 172 180 179 182 181 178 177 186 187 188 184 183 185 191 192 194
+ 190 189 193 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29
+ 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55
+ 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 198 197 196 195 71 72 73 74 75
+ 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119
+ 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 206 203 201 208
+ 202 205 199 207 200 204 210 213 214 212 209 211 219 220 218 217 215 216 223
+ 224 222 225 221 226 229 230 227 228 231 232 237 238 235 236 234 233 241 244
+ 243 242 240 239 247 245 248 246 250 249 251 256 252 255 254 253 262 261 258
+ 260 259 257 265 266 custom_sram_1r1w_32_256_freepdk45_bitcell_array
* cell instance $4 r0 *1 1.175,97.175
X$4 264 263 265 266 custom_sram_1r1w_32_256_freepdk45_dummy_array
.ENDS custom_sram_1r1w_32_256_freepdk45_replica_bitcell_array

* cell custom_sram_1r1w_32_256_freepdk45_pinv
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.1975 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=2.9U AS=0.328425P AD=0.328425P PS=7.575U
+ PD=7.575U
* device instance $21 r0 *1 0.2325,1.1535 PMOS_VTG
M$21 3 1 2 3 PMOS_VTG L=0.05U W=8.65U AS=0.9796125P AD=0.9796125P PS=13.6125U
+ PD=13.6125U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv

* cell custom_sram_1r1w_32_256_freepdk45_pinv_3
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_3 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.17 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.09U AS=0.011475P AD=0.011475P PS=0.435U
+ PD=0.435U
* device instance $2 r0 *1 0.2325,2.21 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_3

* cell custom_sram_1r1w_32_256_freepdk45_pinv_1
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_1 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.185 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.36U AS=0.0423P AD=0.0423P PS=1.185U PD=1.185U
* device instance $4 r0 *1 0.2325,1.19 PMOS_VTG
M$4 3 1 2 3 PMOS_VTG L=0.05U W=1.08U AS=0.1269P AD=0.1269P PS=2.145U PD=2.145U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_1

* cell custom_sram_1r1w_32_256_freepdk45_pnand2
* pin A
* pin B
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pnand2 1 2 3 4 5
* net 1 A
* net 2 B
* net 3 Z
* net 4 vdd
* net 5 gnd
* device instance $1 r0 *1 0.2325,1.235 PMOS_VTG
M$1 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,1.235 PMOS_VTG
M$2 3 2 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.2325,0.215 NMOS_VTG
M$3 5 1 6 5 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $4 r0 *1 0.4475,0.215 NMOS_VTG
M$4 6 2 3 5 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS custom_sram_1r1w_32_256_freepdk45_pnand2

* cell custom_sram_1r1w_32_256_freepdk45_pinv_0
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_pinv_0 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.17 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.09U AS=0.011475P AD=0.011475P PS=0.435U
+ PD=0.435U
* device instance $2 r0 *1 0.2325,1.235 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS custom_sram_1r1w_32_256_freepdk45_pinv_0

* cell custom_sram_1r1w_32_256_freepdk45_replica_column_0
* pin wl_0_0
* pin wl_1_0
* pin wl_1_1
* pin wl_0_1
* pin wl_0_2
* pin wl_1_2
* pin wl_1_3
* pin wl_0_3
* pin wl_0_4
* pin wl_1_4
* pin wl_1_5
* pin wl_0_5
* pin wl_0_6
* pin wl_1_6
* pin wl_1_7
* pin wl_0_7
* pin wl_0_8
* pin wl_1_8
* pin wl_1_9
* pin wl_0_9
* pin wl_0_10
* pin wl_1_10
* pin wl_1_11
* pin wl_0_11
* pin wl_0_12
* pin wl_1_12
* pin wl_1_13
* pin wl_0_13
* pin wl_0_14
* pin wl_1_14
* pin wl_1_15
* pin wl_0_15
* pin wl_0_16
* pin wl_1_16
* pin wl_1_17
* pin wl_0_17
* pin wl_0_18
* pin wl_1_18
* pin wl_1_19
* pin wl_0_19
* pin wl_0_20
* pin wl_1_20
* pin wl_1_21
* pin wl_0_21
* pin wl_0_22
* pin wl_1_22
* pin wl_1_23
* pin wl_0_23
* pin wl_0_24
* pin wl_1_24
* pin wl_1_25
* pin wl_0_25
* pin wl_0_26
* pin wl_1_26
* pin wl_1_27
* pin wl_0_27
* pin wl_0_28
* pin wl_1_28
* pin wl_1_29
* pin wl_0_29
* pin wl_0_30
* pin wl_1_30
* pin wl_1_31
* pin wl_0_31
* pin bl_0_0
* pin bl_1_0
* pin wl_0_32
* pin wl_1_32
* pin br_1_0
* pin br_0_0
* pin wl_1_33
* pin wl_0_33
* pin wl_0_34
* pin wl_1_34
* pin wl_1_35
* pin wl_0_35
* pin wl_0_36
* pin wl_1_36
* pin wl_1_37
* pin wl_0_37
* pin wl_0_38
* pin wl_1_38
* pin wl_1_39
* pin wl_0_39
* pin wl_0_40
* pin wl_1_40
* pin wl_1_41
* pin wl_0_41
* pin wl_0_42
* pin wl_1_42
* pin wl_1_43
* pin wl_0_43
* pin wl_0_44
* pin wl_1_44
* pin wl_1_45
* pin wl_0_45
* pin wl_0_46
* pin wl_1_46
* pin wl_1_47
* pin wl_0_47
* pin wl_0_48
* pin wl_1_48
* pin wl_1_49
* pin wl_0_49
* pin wl_0_50
* pin wl_1_50
* pin wl_1_51
* pin wl_0_51
* pin wl_0_52
* pin wl_1_52
* pin wl_1_53
* pin wl_0_53
* pin wl_0_54
* pin wl_1_54
* pin wl_1_55
* pin wl_0_55
* pin wl_0_56
* pin wl_1_56
* pin wl_1_57
* pin wl_0_57
* pin wl_0_58
* pin wl_1_58
* pin wl_1_59
* pin wl_0_59
* pin wl_0_60
* pin wl_1_60
* pin wl_1_61
* pin wl_0_61
* pin wl_0_62
* pin wl_1_62
* pin wl_1_63
* pin wl_0_63
* pin wl_0_64
* pin wl_1_64
* pin wl_1_65
* pin wl_0_65
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_replica_column_0 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36
+ 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129
+ 130 131 132 133 134 135 136 137 138
* net 1 wl_0_0
* net 2 wl_1_0
* net 3 wl_1_1
* net 4 wl_0_1
* net 5 wl_0_2
* net 6 wl_1_2
* net 7 wl_1_3
* net 8 wl_0_3
* net 9 wl_0_4
* net 10 wl_1_4
* net 11 wl_1_5
* net 12 wl_0_5
* net 13 wl_0_6
* net 14 wl_1_6
* net 15 wl_1_7
* net 16 wl_0_7
* net 17 wl_0_8
* net 18 wl_1_8
* net 19 wl_1_9
* net 20 wl_0_9
* net 21 wl_0_10
* net 22 wl_1_10
* net 23 wl_1_11
* net 24 wl_0_11
* net 25 wl_0_12
* net 26 wl_1_12
* net 27 wl_1_13
* net 28 wl_0_13
* net 29 wl_0_14
* net 30 wl_1_14
* net 31 wl_1_15
* net 32 wl_0_15
* net 33 wl_0_16
* net 34 wl_1_16
* net 35 wl_1_17
* net 36 wl_0_17
* net 37 wl_0_18
* net 38 wl_1_18
* net 39 wl_1_19
* net 40 wl_0_19
* net 41 wl_0_20
* net 42 wl_1_20
* net 43 wl_1_21
* net 44 wl_0_21
* net 45 wl_0_22
* net 46 wl_1_22
* net 47 wl_1_23
* net 48 wl_0_23
* net 49 wl_0_24
* net 50 wl_1_24
* net 51 wl_1_25
* net 52 wl_0_25
* net 53 wl_0_26
* net 54 wl_1_26
* net 55 wl_1_27
* net 56 wl_0_27
* net 57 wl_0_28
* net 58 wl_1_28
* net 59 wl_1_29
* net 60 wl_0_29
* net 61 wl_0_30
* net 62 wl_1_30
* net 63 wl_1_31
* net 64 wl_0_31
* net 65 bl_0_0
* net 66 bl_1_0
* net 67 wl_0_32
* net 68 wl_1_32
* net 69 br_1_0
* net 70 br_0_0
* net 71 wl_1_33
* net 72 wl_0_33
* net 73 wl_0_34
* net 74 wl_1_34
* net 75 wl_1_35
* net 76 wl_0_35
* net 77 wl_0_36
* net 78 wl_1_36
* net 79 wl_1_37
* net 80 wl_0_37
* net 81 wl_0_38
* net 82 wl_1_38
* net 83 wl_1_39
* net 84 wl_0_39
* net 85 wl_0_40
* net 86 wl_1_40
* net 87 wl_1_41
* net 88 wl_0_41
* net 89 wl_0_42
* net 90 wl_1_42
* net 91 wl_1_43
* net 92 wl_0_43
* net 93 wl_0_44
* net 94 wl_1_44
* net 95 wl_1_45
* net 96 wl_0_45
* net 97 wl_0_46
* net 98 wl_1_46
* net 99 wl_1_47
* net 100 wl_0_47
* net 101 wl_0_48
* net 102 wl_1_48
* net 103 wl_1_49
* net 104 wl_0_49
* net 105 wl_0_50
* net 106 wl_1_50
* net 107 wl_1_51
* net 108 wl_0_51
* net 109 wl_0_52
* net 110 wl_1_52
* net 111 wl_1_53
* net 112 wl_0_53
* net 113 wl_0_54
* net 114 wl_1_54
* net 115 wl_1_55
* net 116 wl_0_55
* net 117 wl_0_56
* net 118 wl_1_56
* net 119 wl_1_57
* net 120 wl_0_57
* net 121 wl_0_58
* net 122 wl_1_58
* net 123 wl_1_59
* net 124 wl_0_59
* net 125 wl_0_60
* net 126 wl_1_60
* net 127 wl_1_61
* net 128 wl_0_61
* net 129 wl_0_62
* net 130 wl_1_62
* net 131 wl_1_63
* net 132 wl_0_63
* net 133 wl_0_64
* net 134 wl_1_64
* net 135 wl_1_65
* net 136 wl_0_65
* net 137 vdd
* net 138 gnd
* cell instance $1 m0 *1 0,1.495
X$1 2 1 137 138 dummy_cell_2rw
* cell instance $2 r0 *1 0,1.495
X$2 65 66 69 3 70 4 137 138 replica_cell_2rw
* cell instance $3 m0 *1 0,4.485
X$3 65 66 69 6 70 5 137 138 replica_cell_2rw
* cell instance $4 r0 *1 0,4.485
X$4 65 66 69 7 70 8 137 138 replica_cell_2rw
* cell instance $5 m0 *1 0,7.475
X$5 65 66 69 10 70 9 137 138 replica_cell_2rw
* cell instance $6 r0 *1 0,7.475
X$6 65 66 69 11 70 12 137 138 replica_cell_2rw
* cell instance $7 m0 *1 0,10.465
X$7 65 66 69 14 70 13 137 138 replica_cell_2rw
* cell instance $8 r0 *1 0,10.465
X$8 65 66 69 15 70 16 137 138 replica_cell_2rw
* cell instance $9 m0 *1 0,13.455
X$9 65 66 69 18 70 17 137 138 replica_cell_2rw
* cell instance $10 r0 *1 0,13.455
X$10 65 66 69 19 70 20 137 138 replica_cell_2rw
* cell instance $11 m0 *1 0,16.445
X$11 65 66 69 22 70 21 137 138 replica_cell_2rw
* cell instance $12 r0 *1 0,16.445
X$12 65 66 69 23 70 24 137 138 replica_cell_2rw
* cell instance $13 m0 *1 0,19.435
X$13 65 66 69 26 70 25 137 138 replica_cell_2rw
* cell instance $14 r0 *1 0,19.435
X$14 65 66 69 27 70 28 137 138 replica_cell_2rw
* cell instance $15 m0 *1 0,22.425
X$15 65 66 69 30 70 29 137 138 replica_cell_2rw
* cell instance $16 r0 *1 0,22.425
X$16 65 66 69 31 70 32 137 138 replica_cell_2rw
* cell instance $17 m0 *1 0,25.415
X$17 65 66 69 34 70 33 137 138 replica_cell_2rw
* cell instance $18 r0 *1 0,25.415
X$18 65 66 69 35 70 36 137 138 replica_cell_2rw
* cell instance $19 m0 *1 0,28.405
X$19 65 66 69 38 70 37 137 138 replica_cell_2rw
* cell instance $20 r0 *1 0,28.405
X$20 65 66 69 39 70 40 137 138 replica_cell_2rw
* cell instance $21 m0 *1 0,31.395
X$21 65 66 69 42 70 41 137 138 replica_cell_2rw
* cell instance $22 r0 *1 0,31.395
X$22 65 66 69 43 70 44 137 138 replica_cell_2rw
* cell instance $23 m0 *1 0,34.385
X$23 65 66 69 46 70 45 137 138 replica_cell_2rw
* cell instance $24 r0 *1 0,34.385
X$24 65 66 69 47 70 48 137 138 replica_cell_2rw
* cell instance $25 m0 *1 0,37.375
X$25 65 66 69 50 70 49 137 138 replica_cell_2rw
* cell instance $26 r0 *1 0,37.375
X$26 65 66 69 51 70 52 137 138 replica_cell_2rw
* cell instance $27 m0 *1 0,40.365
X$27 65 66 69 54 70 53 137 138 replica_cell_2rw
* cell instance $28 r0 *1 0,40.365
X$28 65 66 69 55 70 56 137 138 replica_cell_2rw
* cell instance $29 m0 *1 0,43.355
X$29 65 66 69 58 70 57 137 138 replica_cell_2rw
* cell instance $30 r0 *1 0,43.355
X$30 65 66 69 59 70 60 137 138 replica_cell_2rw
* cell instance $31 m0 *1 0,46.345
X$31 65 66 69 62 70 61 137 138 replica_cell_2rw
* cell instance $32 r0 *1 0,46.345
X$32 65 66 69 63 70 64 137 138 replica_cell_2rw
* cell instance $33 m0 *1 0,49.335
X$33 65 66 69 68 70 67 137 138 replica_cell_2rw
* cell instance $34 r0 *1 0,49.335
X$34 65 66 69 71 70 72 137 138 replica_cell_2rw
* cell instance $35 m0 *1 0,52.325
X$35 65 66 69 74 70 73 137 138 replica_cell_2rw
* cell instance $36 r0 *1 0,52.325
X$36 65 66 69 75 70 76 137 138 replica_cell_2rw
* cell instance $37 m0 *1 0,55.315
X$37 65 66 69 78 70 77 137 138 replica_cell_2rw
* cell instance $38 r0 *1 0,55.315
X$38 65 66 69 79 70 80 137 138 replica_cell_2rw
* cell instance $39 m0 *1 0,58.305
X$39 65 66 69 82 70 81 137 138 replica_cell_2rw
* cell instance $40 r0 *1 0,58.305
X$40 65 66 69 83 70 84 137 138 replica_cell_2rw
* cell instance $41 m0 *1 0,61.295
X$41 65 66 69 86 70 85 137 138 replica_cell_2rw
* cell instance $42 r0 *1 0,61.295
X$42 65 66 69 87 70 88 137 138 replica_cell_2rw
* cell instance $43 m0 *1 0,64.285
X$43 65 66 69 90 70 89 137 138 replica_cell_2rw
* cell instance $44 r0 *1 0,64.285
X$44 65 66 69 91 70 92 137 138 replica_cell_2rw
* cell instance $45 m0 *1 0,67.275
X$45 65 66 69 94 70 93 137 138 replica_cell_2rw
* cell instance $46 r0 *1 0,67.275
X$46 65 66 69 95 70 96 137 138 replica_cell_2rw
* cell instance $47 m0 *1 0,70.265
X$47 65 66 69 98 70 97 137 138 replica_cell_2rw
* cell instance $48 r0 *1 0,70.265
X$48 65 66 69 99 70 100 137 138 replica_cell_2rw
* cell instance $49 m0 *1 0,73.255
X$49 65 66 69 102 70 101 137 138 replica_cell_2rw
* cell instance $50 r0 *1 0,73.255
X$50 65 66 69 103 70 104 137 138 replica_cell_2rw
* cell instance $51 m0 *1 0,76.245
X$51 65 66 69 106 70 105 137 138 replica_cell_2rw
* cell instance $52 r0 *1 0,76.245
X$52 65 66 69 107 70 108 137 138 replica_cell_2rw
* cell instance $53 m0 *1 0,79.235
X$53 65 66 69 110 70 109 137 138 replica_cell_2rw
* cell instance $54 r0 *1 0,79.235
X$54 65 66 69 111 70 112 137 138 replica_cell_2rw
* cell instance $55 m0 *1 0,82.225
X$55 65 66 69 114 70 113 137 138 replica_cell_2rw
* cell instance $56 r0 *1 0,82.225
X$56 65 66 69 115 70 116 137 138 replica_cell_2rw
* cell instance $57 m0 *1 0,85.215
X$57 65 66 69 118 70 117 137 138 replica_cell_2rw
* cell instance $58 r0 *1 0,85.215
X$58 65 66 69 119 70 120 137 138 replica_cell_2rw
* cell instance $59 m0 *1 0,88.205
X$59 65 66 69 122 70 121 137 138 replica_cell_2rw
* cell instance $60 r0 *1 0,88.205
X$60 65 66 69 123 70 124 137 138 replica_cell_2rw
* cell instance $61 m0 *1 0,91.195
X$61 65 66 69 126 70 125 137 138 replica_cell_2rw
* cell instance $62 r0 *1 0,91.195
X$62 65 66 69 127 70 128 137 138 replica_cell_2rw
* cell instance $63 m0 *1 0,94.185
X$63 65 66 69 130 70 129 137 138 replica_cell_2rw
* cell instance $64 r0 *1 0,94.185
X$64 65 66 69 131 70 132 137 138 replica_cell_2rw
* cell instance $65 m0 *1 0,97.175
X$65 65 66 69 134 70 133 137 138 replica_cell_2rw
* cell instance $66 r0 *1 0,97.175
X$66 65 66 69 135 70 136 137 138 replica_cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_replica_column_0

* cell custom_sram_1r1w_32_256_freepdk45_dummy_array_4
* pin wl_0_0
* pin wl_1_0
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_dummy_array_4 1 2 3 4
* net 1 wl_0_0
* net 2 wl_1_0
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 dummy_cell_2rw
* cell instance $2 r0 *1 1.175,0
X$2 2 1 3 4 dummy_cell_2rw
* cell instance $3 r0 *1 2.35,0
X$3 2 1 3 4 dummy_cell_2rw
* cell instance $4 r0 *1 3.525,0
X$4 2 1 3 4 dummy_cell_2rw
* cell instance $5 r0 *1 4.7,0
X$5 2 1 3 4 dummy_cell_2rw
* cell instance $6 r0 *1 5.875,0
X$6 2 1 3 4 dummy_cell_2rw
* cell instance $7 r0 *1 7.05,0
X$7 2 1 3 4 dummy_cell_2rw
* cell instance $8 r0 *1 8.225,0
X$8 2 1 3 4 dummy_cell_2rw
* cell instance $9 r0 *1 9.4,0
X$9 2 1 3 4 dummy_cell_2rw
* cell instance $10 r0 *1 10.575,0
X$10 2 1 3 4 dummy_cell_2rw
* cell instance $11 r0 *1 11.75,0
X$11 2 1 3 4 dummy_cell_2rw
* cell instance $12 r0 *1 12.925,0
X$12 2 1 3 4 dummy_cell_2rw
* cell instance $13 r0 *1 14.1,0
X$13 2 1 3 4 dummy_cell_2rw
* cell instance $14 r0 *1 15.275,0
X$14 2 1 3 4 dummy_cell_2rw
* cell instance $15 r0 *1 16.45,0
X$15 2 1 3 4 dummy_cell_2rw
* cell instance $16 r0 *1 17.625,0
X$16 2 1 3 4 dummy_cell_2rw
* cell instance $17 r0 *1 18.8,0
X$17 2 1 3 4 dummy_cell_2rw
* cell instance $18 r0 *1 19.975,0
X$18 2 1 3 4 dummy_cell_2rw
* cell instance $19 r0 *1 21.15,0
X$19 2 1 3 4 dummy_cell_2rw
* cell instance $20 r0 *1 22.325,0
X$20 2 1 3 4 dummy_cell_2rw
* cell instance $21 r0 *1 23.5,0
X$21 2 1 3 4 dummy_cell_2rw
* cell instance $22 r0 *1 24.675,0
X$22 2 1 3 4 dummy_cell_2rw
* cell instance $23 r0 *1 25.85,0
X$23 2 1 3 4 dummy_cell_2rw
* cell instance $24 r0 *1 27.025,0
X$24 2 1 3 4 dummy_cell_2rw
* cell instance $25 r0 *1 28.2,0
X$25 2 1 3 4 dummy_cell_2rw
* cell instance $26 r0 *1 29.375,0
X$26 2 1 3 4 dummy_cell_2rw
* cell instance $27 r0 *1 30.55,0
X$27 2 1 3 4 dummy_cell_2rw
* cell instance $28 r0 *1 31.725,0
X$28 2 1 3 4 dummy_cell_2rw
* cell instance $29 r0 *1 32.9,0
X$29 2 1 3 4 dummy_cell_2rw
* cell instance $30 r0 *1 34.075,0
X$30 2 1 3 4 dummy_cell_2rw
* cell instance $31 r0 *1 35.25,0
X$31 2 1 3 4 dummy_cell_2rw
* cell instance $32 r0 *1 36.425,0
X$32 2 1 3 4 dummy_cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_dummy_array_4

* cell custom_sram_1r1w_32_256_freepdk45_bitcell_array_0
* pin wl_0_2
* pin wl_1_2
* pin wl_0_1
* pin wl_1_1
* pin wl_0_0
* pin wl_1_0
* pin wl_1_4
* pin wl_0_5
* pin wl_1_5
* pin wl_0_4
* pin wl_1_3
* pin wl_0_3
* pin wl_1_7
* pin wl_0_7
* pin wl_0_8
* pin wl_1_8
* pin wl_1_6
* pin wl_0_6
* pin wl_0_10
* pin wl_1_10
* pin wl_1_11
* pin wl_0_11
* pin wl_0_9
* pin wl_1_9
* pin wl_0_14
* pin wl_1_13
* pin wl_1_12
* pin wl_1_14
* pin wl_0_13
* pin wl_0_12
* pin wl_1_16
* pin wl_0_17
* pin wl_0_16
* pin wl_1_17
* pin wl_1_15
* pin wl_0_15
* pin wl_1_20
* pin wl_0_20
* pin wl_0_18
* pin wl_0_19
* pin wl_1_19
* pin wl_1_18
* pin wl_0_22
* pin wl_1_22
* pin wl_1_23
* pin wl_0_23
* pin wl_0_21
* pin wl_1_21
* pin wl_0_25
* pin wl_0_26
* pin wl_1_26
* pin wl_0_24
* pin wl_1_24
* pin wl_1_25
* pin wl_0_28
* pin wl_1_28
* pin wl_0_29
* pin wl_0_27
* pin wl_1_27
* pin wl_1_29
* pin bl_0_0
* pin bl_1_0
* pin br_1_0
* pin br_0_0
* pin bl_0_1
* pin bl_1_1
* pin br_1_1
* pin br_0_1
* pin bl_0_2
* pin bl_1_2
* pin br_1_2
* pin br_0_2
* pin bl_0_3
* pin bl_1_3
* pin br_1_3
* pin br_0_3
* pin bl_0_4
* pin bl_1_4
* pin br_1_4
* pin br_0_4
* pin bl_0_5
* pin bl_1_5
* pin br_1_5
* pin br_0_5
* pin bl_0_6
* pin bl_1_6
* pin br_1_6
* pin br_0_6
* pin bl_0_7
* pin bl_1_7
* pin br_1_7
* pin br_0_7
* pin bl_0_8
* pin bl_1_8
* pin br_1_8
* pin br_0_8
* pin bl_0_9
* pin bl_1_9
* pin br_1_9
* pin br_0_9
* pin bl_0_10
* pin bl_1_10
* pin br_1_10
* pin br_0_10
* pin bl_0_11
* pin bl_1_11
* pin br_1_11
* pin br_0_11
* pin bl_0_12
* pin bl_1_12
* pin br_1_12
* pin br_0_12
* pin bl_0_13
* pin bl_1_13
* pin br_1_13
* pin br_0_13
* pin bl_0_14
* pin bl_1_14
* pin br_1_14
* pin br_0_14
* pin bl_0_15
* pin bl_1_15
* pin br_1_15
* pin br_0_15
* pin wl_0_31
* pin wl_1_31
* pin wl_1_30
* pin wl_0_30
* pin bl_0_16
* pin bl_1_16
* pin br_1_16
* pin br_0_16
* pin bl_0_17
* pin bl_1_17
* pin br_1_17
* pin br_0_17
* pin bl_0_18
* pin bl_1_18
* pin br_1_18
* pin br_0_18
* pin bl_0_19
* pin bl_1_19
* pin br_1_19
* pin br_0_19
* pin bl_0_20
* pin bl_1_20
* pin br_1_20
* pin br_0_20
* pin bl_0_21
* pin bl_1_21
* pin br_1_21
* pin br_0_21
* pin bl_0_22
* pin bl_1_22
* pin br_1_22
* pin br_0_22
* pin bl_0_23
* pin bl_1_23
* pin br_1_23
* pin br_0_23
* pin bl_0_24
* pin bl_1_24
* pin br_1_24
* pin br_0_24
* pin bl_0_25
* pin bl_1_25
* pin br_1_25
* pin br_0_25
* pin bl_0_26
* pin bl_1_26
* pin br_1_26
* pin br_0_26
* pin bl_0_27
* pin bl_1_27
* pin br_1_27
* pin br_0_27
* pin bl_0_28
* pin bl_1_28
* pin br_1_28
* pin br_0_28
* pin bl_0_29
* pin bl_1_29
* pin br_1_29
* pin br_0_29
* pin bl_0_30
* pin bl_1_30
* pin br_1_30
* pin br_0_30
* pin bl_0_31
* pin bl_1_31
* pin br_1_31
* pin br_0_31
* pin wl_0_35
* pin wl_0_34
* pin wl_1_33
* pin wl_1_36
* pin wl_0_33
* pin wl_1_35
* pin wl_1_32
* pin wl_0_36
* pin wl_0_32
* pin wl_1_34
* pin wl_1_37
* pin wl_0_39
* pin wl_1_39
* pin wl_1_38
* pin wl_0_37
* pin wl_0_38
* pin wl_0_42
* pin wl_1_42
* pin wl_0_41
* pin wl_1_41
* pin wl_0_40
* pin wl_1_40
* pin wl_0_44
* pin wl_1_44
* pin wl_0_43
* pin wl_1_45
* pin wl_1_43
* pin wl_0_45
* pin wl_1_47
* pin wl_0_47
* pin wl_0_46
* pin wl_1_46
* pin wl_0_48
* pin wl_1_48
* pin wl_1_51
* pin wl_0_51
* pin wl_0_50
* pin wl_1_50
* pin wl_1_49
* pin wl_0_49
* pin wl_1_53
* pin wl_0_54
* pin wl_1_54
* pin wl_0_53
* pin wl_1_52
* pin wl_0_52
* pin wl_1_56
* pin wl_1_55
* pin wl_0_56
* pin wl_0_55
* pin wl_0_57
* pin wl_1_57
* pin wl_1_58
* pin wl_1_60
* pin wl_0_58
* pin wl_0_60
* pin wl_0_59
* pin wl_1_59
* pin wl_1_63
* pin wl_0_63
* pin wl_1_61
* pin wl_0_62
* pin wl_1_62
* pin wl_0_61
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_bitcell_array_0 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36
+ 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129
+ 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148
+ 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167
+ 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186
+ 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205
+ 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224
+ 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243
+ 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258
* net 1 wl_0_2
* net 2 wl_1_2
* net 3 wl_0_1
* net 4 wl_1_1
* net 5 wl_0_0
* net 6 wl_1_0
* net 7 wl_1_4
* net 8 wl_0_5
* net 9 wl_1_5
* net 10 wl_0_4
* net 11 wl_1_3
* net 12 wl_0_3
* net 13 wl_1_7
* net 14 wl_0_7
* net 15 wl_0_8
* net 16 wl_1_8
* net 17 wl_1_6
* net 18 wl_0_6
* net 19 wl_0_10
* net 20 wl_1_10
* net 21 wl_1_11
* net 22 wl_0_11
* net 23 wl_0_9
* net 24 wl_1_9
* net 25 wl_0_14
* net 26 wl_1_13
* net 27 wl_1_12
* net 28 wl_1_14
* net 29 wl_0_13
* net 30 wl_0_12
* net 31 wl_1_16
* net 32 wl_0_17
* net 33 wl_0_16
* net 34 wl_1_17
* net 35 wl_1_15
* net 36 wl_0_15
* net 37 wl_1_20
* net 38 wl_0_20
* net 39 wl_0_18
* net 40 wl_0_19
* net 41 wl_1_19
* net 42 wl_1_18
* net 43 wl_0_22
* net 44 wl_1_22
* net 45 wl_1_23
* net 46 wl_0_23
* net 47 wl_0_21
* net 48 wl_1_21
* net 49 wl_0_25
* net 50 wl_0_26
* net 51 wl_1_26
* net 52 wl_0_24
* net 53 wl_1_24
* net 54 wl_1_25
* net 55 wl_0_28
* net 56 wl_1_28
* net 57 wl_0_29
* net 58 wl_0_27
* net 59 wl_1_27
* net 60 wl_1_29
* net 61 bl_0_0
* net 62 bl_1_0
* net 63 br_1_0
* net 64 br_0_0
* net 65 bl_0_1
* net 66 bl_1_1
* net 67 br_1_1
* net 68 br_0_1
* net 69 bl_0_2
* net 70 bl_1_2
* net 71 br_1_2
* net 72 br_0_2
* net 73 bl_0_3
* net 74 bl_1_3
* net 75 br_1_3
* net 76 br_0_3
* net 77 bl_0_4
* net 78 bl_1_4
* net 79 br_1_4
* net 80 br_0_4
* net 81 bl_0_5
* net 82 bl_1_5
* net 83 br_1_5
* net 84 br_0_5
* net 85 bl_0_6
* net 86 bl_1_6
* net 87 br_1_6
* net 88 br_0_6
* net 89 bl_0_7
* net 90 bl_1_7
* net 91 br_1_7
* net 92 br_0_7
* net 93 bl_0_8
* net 94 bl_1_8
* net 95 br_1_8
* net 96 br_0_8
* net 97 bl_0_9
* net 98 bl_1_9
* net 99 br_1_9
* net 100 br_0_9
* net 101 bl_0_10
* net 102 bl_1_10
* net 103 br_1_10
* net 104 br_0_10
* net 105 bl_0_11
* net 106 bl_1_11
* net 107 br_1_11
* net 108 br_0_11
* net 109 bl_0_12
* net 110 bl_1_12
* net 111 br_1_12
* net 112 br_0_12
* net 113 bl_0_13
* net 114 bl_1_13
* net 115 br_1_13
* net 116 br_0_13
* net 117 bl_0_14
* net 118 bl_1_14
* net 119 br_1_14
* net 120 br_0_14
* net 121 bl_0_15
* net 122 bl_1_15
* net 123 br_1_15
* net 124 br_0_15
* net 125 wl_0_31
* net 126 wl_1_31
* net 127 wl_1_30
* net 128 wl_0_30
* net 129 bl_0_16
* net 130 bl_1_16
* net 131 br_1_16
* net 132 br_0_16
* net 133 bl_0_17
* net 134 bl_1_17
* net 135 br_1_17
* net 136 br_0_17
* net 137 bl_0_18
* net 138 bl_1_18
* net 139 br_1_18
* net 140 br_0_18
* net 141 bl_0_19
* net 142 bl_1_19
* net 143 br_1_19
* net 144 br_0_19
* net 145 bl_0_20
* net 146 bl_1_20
* net 147 br_1_20
* net 148 br_0_20
* net 149 bl_0_21
* net 150 bl_1_21
* net 151 br_1_21
* net 152 br_0_21
* net 153 bl_0_22
* net 154 bl_1_22
* net 155 br_1_22
* net 156 br_0_22
* net 157 bl_0_23
* net 158 bl_1_23
* net 159 br_1_23
* net 160 br_0_23
* net 161 bl_0_24
* net 162 bl_1_24
* net 163 br_1_24
* net 164 br_0_24
* net 165 bl_0_25
* net 166 bl_1_25
* net 167 br_1_25
* net 168 br_0_25
* net 169 bl_0_26
* net 170 bl_1_26
* net 171 br_1_26
* net 172 br_0_26
* net 173 bl_0_27
* net 174 bl_1_27
* net 175 br_1_27
* net 176 br_0_27
* net 177 bl_0_28
* net 178 bl_1_28
* net 179 br_1_28
* net 180 br_0_28
* net 181 bl_0_29
* net 182 bl_1_29
* net 183 br_1_29
* net 184 br_0_29
* net 185 bl_0_30
* net 186 bl_1_30
* net 187 br_1_30
* net 188 br_0_30
* net 189 bl_0_31
* net 190 bl_1_31
* net 191 br_1_31
* net 192 br_0_31
* net 193 wl_0_35
* net 194 wl_0_34
* net 195 wl_1_33
* net 196 wl_1_36
* net 197 wl_0_33
* net 198 wl_1_35
* net 199 wl_1_32
* net 200 wl_0_36
* net 201 wl_0_32
* net 202 wl_1_34
* net 203 wl_1_37
* net 204 wl_0_39
* net 205 wl_1_39
* net 206 wl_1_38
* net 207 wl_0_37
* net 208 wl_0_38
* net 209 wl_0_42
* net 210 wl_1_42
* net 211 wl_0_41
* net 212 wl_1_41
* net 213 wl_0_40
* net 214 wl_1_40
* net 215 wl_0_44
* net 216 wl_1_44
* net 217 wl_0_43
* net 218 wl_1_45
* net 219 wl_1_43
* net 220 wl_0_45
* net 221 wl_1_47
* net 222 wl_0_47
* net 223 wl_0_46
* net 224 wl_1_46
* net 225 wl_0_48
* net 226 wl_1_48
* net 227 wl_1_51
* net 228 wl_0_51
* net 229 wl_0_50
* net 230 wl_1_50
* net 231 wl_1_49
* net 232 wl_0_49
* net 233 wl_1_53
* net 234 wl_0_54
* net 235 wl_1_54
* net 236 wl_0_53
* net 237 wl_1_52
* net 238 wl_0_52
* net 239 wl_1_56
* net 240 wl_1_55
* net 241 wl_0_56
* net 242 wl_0_55
* net 243 wl_0_57
* net 244 wl_1_57
* net 245 wl_1_58
* net 246 wl_1_60
* net 247 wl_0_58
* net 248 wl_0_60
* net 249 wl_0_59
* net 250 wl_1_59
* net 251 wl_1_63
* net 252 wl_0_63
* net 253 wl_1_61
* net 254 wl_0_62
* net 255 wl_1_62
* net 256 wl_0_61
* net 257 vdd
* net 258 gnd
* cell instance $1 r0 *1 1.175,2.99
X$1 65 66 67 2 68 1 257 258 cell_2rw
* cell instance $2 r0 *1 0,2.99
X$2 61 62 63 2 64 1 257 258 cell_2rw
* cell instance $3 r0 *1 2.35,2.99
X$3 69 70 71 2 72 1 257 258 cell_2rw
* cell instance $4 r0 *1 3.525,2.99
X$4 73 74 75 2 76 1 257 258 cell_2rw
* cell instance $5 r0 *1 4.7,2.99
X$5 77 78 79 2 80 1 257 258 cell_2rw
* cell instance $6 r0 *1 5.875,2.99
X$6 81 82 83 2 84 1 257 258 cell_2rw
* cell instance $7 r0 *1 7.05,2.99
X$7 85 86 87 2 88 1 257 258 cell_2rw
* cell instance $8 r0 *1 8.225,2.99
X$8 89 90 91 2 92 1 257 258 cell_2rw
* cell instance $9 r0 *1 9.4,2.99
X$9 93 94 95 2 96 1 257 258 cell_2rw
* cell instance $10 r0 *1 10.575,2.99
X$10 97 98 99 2 100 1 257 258 cell_2rw
* cell instance $11 r0 *1 11.75,2.99
X$11 101 102 103 2 104 1 257 258 cell_2rw
* cell instance $12 r0 *1 12.925,2.99
X$12 105 106 107 2 108 1 257 258 cell_2rw
* cell instance $13 r0 *1 14.1,2.99
X$13 109 110 111 2 112 1 257 258 cell_2rw
* cell instance $14 r0 *1 15.275,2.99
X$14 113 114 115 2 116 1 257 258 cell_2rw
* cell instance $15 r0 *1 16.45,2.99
X$15 117 118 119 2 120 1 257 258 cell_2rw
* cell instance $16 r0 *1 17.625,2.99
X$16 121 122 123 2 124 1 257 258 cell_2rw
* cell instance $17 r0 *1 18.8,2.99
X$17 129 130 131 2 132 1 257 258 cell_2rw
* cell instance $18 r0 *1 19.975,2.99
X$18 133 134 135 2 136 1 257 258 cell_2rw
* cell instance $19 r0 *1 21.15,2.99
X$19 137 138 139 2 140 1 257 258 cell_2rw
* cell instance $20 r0 *1 22.325,2.99
X$20 141 142 143 2 144 1 257 258 cell_2rw
* cell instance $21 r0 *1 23.5,2.99
X$21 145 146 147 2 148 1 257 258 cell_2rw
* cell instance $22 r0 *1 24.675,2.99
X$22 149 150 151 2 152 1 257 258 cell_2rw
* cell instance $23 r0 *1 25.85,2.99
X$23 153 154 155 2 156 1 257 258 cell_2rw
* cell instance $24 r0 *1 27.025,2.99
X$24 157 158 159 2 160 1 257 258 cell_2rw
* cell instance $25 r0 *1 28.2,2.99
X$25 161 162 163 2 164 1 257 258 cell_2rw
* cell instance $26 r0 *1 29.375,2.99
X$26 165 166 167 2 168 1 257 258 cell_2rw
* cell instance $27 r0 *1 30.55,2.99
X$27 169 170 171 2 172 1 257 258 cell_2rw
* cell instance $28 r0 *1 31.725,2.99
X$28 173 174 175 2 176 1 257 258 cell_2rw
* cell instance $29 r0 *1 32.9,2.99
X$29 177 178 179 2 180 1 257 258 cell_2rw
* cell instance $30 r0 *1 34.075,2.99
X$30 181 182 183 2 184 1 257 258 cell_2rw
* cell instance $31 r0 *1 35.25,2.99
X$31 185 186 187 2 188 1 257 258 cell_2rw
* cell instance $32 r0 *1 36.425,2.99
X$32 189 190 191 2 192 1 257 258 cell_2rw
* cell instance $33 m0 *1 1.175,2.99
X$33 65 66 67 4 68 3 257 258 cell_2rw
* cell instance $34 m0 *1 0,2.99
X$34 61 62 63 4 64 3 257 258 cell_2rw
* cell instance $35 m0 *1 2.35,2.99
X$35 69 70 71 4 72 3 257 258 cell_2rw
* cell instance $36 m0 *1 3.525,2.99
X$36 73 74 75 4 76 3 257 258 cell_2rw
* cell instance $37 m0 *1 4.7,2.99
X$37 77 78 79 4 80 3 257 258 cell_2rw
* cell instance $38 m0 *1 5.875,2.99
X$38 81 82 83 4 84 3 257 258 cell_2rw
* cell instance $39 m0 *1 7.05,2.99
X$39 85 86 87 4 88 3 257 258 cell_2rw
* cell instance $40 m0 *1 8.225,2.99
X$40 89 90 91 4 92 3 257 258 cell_2rw
* cell instance $41 m0 *1 9.4,2.99
X$41 93 94 95 4 96 3 257 258 cell_2rw
* cell instance $42 m0 *1 10.575,2.99
X$42 97 98 99 4 100 3 257 258 cell_2rw
* cell instance $43 m0 *1 11.75,2.99
X$43 101 102 103 4 104 3 257 258 cell_2rw
* cell instance $44 m0 *1 12.925,2.99
X$44 105 106 107 4 108 3 257 258 cell_2rw
* cell instance $45 m0 *1 14.1,2.99
X$45 109 110 111 4 112 3 257 258 cell_2rw
* cell instance $46 m0 *1 15.275,2.99
X$46 113 114 115 4 116 3 257 258 cell_2rw
* cell instance $47 m0 *1 16.45,2.99
X$47 117 118 119 4 120 3 257 258 cell_2rw
* cell instance $48 m0 *1 17.625,2.99
X$48 121 122 123 4 124 3 257 258 cell_2rw
* cell instance $49 m0 *1 18.8,2.99
X$49 129 130 131 4 132 3 257 258 cell_2rw
* cell instance $50 m0 *1 19.975,2.99
X$50 133 134 135 4 136 3 257 258 cell_2rw
* cell instance $51 m0 *1 21.15,2.99
X$51 137 138 139 4 140 3 257 258 cell_2rw
* cell instance $52 m0 *1 22.325,2.99
X$52 141 142 143 4 144 3 257 258 cell_2rw
* cell instance $53 m0 *1 23.5,2.99
X$53 145 146 147 4 148 3 257 258 cell_2rw
* cell instance $54 m0 *1 24.675,2.99
X$54 149 150 151 4 152 3 257 258 cell_2rw
* cell instance $55 m0 *1 25.85,2.99
X$55 153 154 155 4 156 3 257 258 cell_2rw
* cell instance $56 m0 *1 27.025,2.99
X$56 157 158 159 4 160 3 257 258 cell_2rw
* cell instance $57 m0 *1 28.2,2.99
X$57 161 162 163 4 164 3 257 258 cell_2rw
* cell instance $58 m0 *1 29.375,2.99
X$58 165 166 167 4 168 3 257 258 cell_2rw
* cell instance $59 m0 *1 30.55,2.99
X$59 169 170 171 4 172 3 257 258 cell_2rw
* cell instance $60 m0 *1 31.725,2.99
X$60 173 174 175 4 176 3 257 258 cell_2rw
* cell instance $61 m0 *1 32.9,2.99
X$61 177 178 179 4 180 3 257 258 cell_2rw
* cell instance $62 m0 *1 34.075,2.99
X$62 181 182 183 4 184 3 257 258 cell_2rw
* cell instance $63 m0 *1 35.25,2.99
X$63 185 186 187 4 188 3 257 258 cell_2rw
* cell instance $64 m0 *1 36.425,2.99
X$64 189 190 191 4 192 3 257 258 cell_2rw
* cell instance $65 r0 *1 0,0
X$65 61 62 63 6 64 5 257 258 cell_2rw
* cell instance $66 r0 *1 1.175,0
X$66 65 66 67 6 68 5 257 258 cell_2rw
* cell instance $67 r0 *1 2.35,0
X$67 69 70 71 6 72 5 257 258 cell_2rw
* cell instance $68 r0 *1 3.525,0
X$68 73 74 75 6 76 5 257 258 cell_2rw
* cell instance $69 r0 *1 4.7,0
X$69 77 78 79 6 80 5 257 258 cell_2rw
* cell instance $70 r0 *1 5.875,0
X$70 81 82 83 6 84 5 257 258 cell_2rw
* cell instance $71 r0 *1 7.05,0
X$71 85 86 87 6 88 5 257 258 cell_2rw
* cell instance $72 r0 *1 8.225,0
X$72 89 90 91 6 92 5 257 258 cell_2rw
* cell instance $73 r0 *1 9.4,0
X$73 93 94 95 6 96 5 257 258 cell_2rw
* cell instance $74 r0 *1 10.575,0
X$74 97 98 99 6 100 5 257 258 cell_2rw
* cell instance $75 r0 *1 11.75,0
X$75 101 102 103 6 104 5 257 258 cell_2rw
* cell instance $76 r0 *1 12.925,0
X$76 105 106 107 6 108 5 257 258 cell_2rw
* cell instance $77 r0 *1 14.1,0
X$77 109 110 111 6 112 5 257 258 cell_2rw
* cell instance $78 r0 *1 15.275,0
X$78 113 114 115 6 116 5 257 258 cell_2rw
* cell instance $79 r0 *1 16.45,0
X$79 117 118 119 6 120 5 257 258 cell_2rw
* cell instance $80 r0 *1 17.625,0
X$80 121 122 123 6 124 5 257 258 cell_2rw
* cell instance $81 r0 *1 18.8,0
X$81 129 130 131 6 132 5 257 258 cell_2rw
* cell instance $82 r0 *1 19.975,0
X$82 133 134 135 6 136 5 257 258 cell_2rw
* cell instance $83 r0 *1 21.15,0
X$83 137 138 139 6 140 5 257 258 cell_2rw
* cell instance $84 r0 *1 22.325,0
X$84 141 142 143 6 144 5 257 258 cell_2rw
* cell instance $85 r0 *1 23.5,0
X$85 145 146 147 6 148 5 257 258 cell_2rw
* cell instance $86 r0 *1 24.675,0
X$86 149 150 151 6 152 5 257 258 cell_2rw
* cell instance $87 r0 *1 25.85,0
X$87 153 154 155 6 156 5 257 258 cell_2rw
* cell instance $88 r0 *1 27.025,0
X$88 157 158 159 6 160 5 257 258 cell_2rw
* cell instance $89 r0 *1 28.2,0
X$89 161 162 163 6 164 5 257 258 cell_2rw
* cell instance $90 r0 *1 29.375,0
X$90 165 166 167 6 168 5 257 258 cell_2rw
* cell instance $91 r0 *1 30.55,0
X$91 169 170 171 6 172 5 257 258 cell_2rw
* cell instance $92 r0 *1 31.725,0
X$92 173 174 175 6 176 5 257 258 cell_2rw
* cell instance $93 r0 *1 32.9,0
X$93 177 178 179 6 180 5 257 258 cell_2rw
* cell instance $94 r0 *1 34.075,0
X$94 181 182 183 6 184 5 257 258 cell_2rw
* cell instance $95 r0 *1 35.25,0
X$95 185 186 187 6 188 5 257 258 cell_2rw
* cell instance $96 r0 *1 36.425,0
X$96 189 190 191 6 192 5 257 258 cell_2rw
* cell instance $97 r0 *1 1.175,5.98
X$97 65 66 67 7 68 10 257 258 cell_2rw
* cell instance $98 r0 *1 0,5.98
X$98 61 62 63 7 64 10 257 258 cell_2rw
* cell instance $99 r0 *1 2.35,5.98
X$99 69 70 71 7 72 10 257 258 cell_2rw
* cell instance $100 r0 *1 3.525,5.98
X$100 73 74 75 7 76 10 257 258 cell_2rw
* cell instance $101 r0 *1 4.7,5.98
X$101 77 78 79 7 80 10 257 258 cell_2rw
* cell instance $102 r0 *1 5.875,5.98
X$102 81 82 83 7 84 10 257 258 cell_2rw
* cell instance $103 r0 *1 7.05,5.98
X$103 85 86 87 7 88 10 257 258 cell_2rw
* cell instance $104 r0 *1 8.225,5.98
X$104 89 90 91 7 92 10 257 258 cell_2rw
* cell instance $105 r0 *1 9.4,5.98
X$105 93 94 95 7 96 10 257 258 cell_2rw
* cell instance $106 r0 *1 10.575,5.98
X$106 97 98 99 7 100 10 257 258 cell_2rw
* cell instance $107 r0 *1 11.75,5.98
X$107 101 102 103 7 104 10 257 258 cell_2rw
* cell instance $108 r0 *1 12.925,5.98
X$108 105 106 107 7 108 10 257 258 cell_2rw
* cell instance $109 r0 *1 14.1,5.98
X$109 109 110 111 7 112 10 257 258 cell_2rw
* cell instance $110 r0 *1 15.275,5.98
X$110 113 114 115 7 116 10 257 258 cell_2rw
* cell instance $111 r0 *1 16.45,5.98
X$111 117 118 119 7 120 10 257 258 cell_2rw
* cell instance $112 r0 *1 17.625,5.98
X$112 121 122 123 7 124 10 257 258 cell_2rw
* cell instance $113 r0 *1 18.8,5.98
X$113 129 130 131 7 132 10 257 258 cell_2rw
* cell instance $114 r0 *1 19.975,5.98
X$114 133 134 135 7 136 10 257 258 cell_2rw
* cell instance $115 r0 *1 21.15,5.98
X$115 137 138 139 7 140 10 257 258 cell_2rw
* cell instance $116 r0 *1 22.325,5.98
X$116 141 142 143 7 144 10 257 258 cell_2rw
* cell instance $117 r0 *1 23.5,5.98
X$117 145 146 147 7 148 10 257 258 cell_2rw
* cell instance $118 r0 *1 24.675,5.98
X$118 149 150 151 7 152 10 257 258 cell_2rw
* cell instance $119 r0 *1 25.85,5.98
X$119 153 154 155 7 156 10 257 258 cell_2rw
* cell instance $120 r0 *1 27.025,5.98
X$120 157 158 159 7 160 10 257 258 cell_2rw
* cell instance $121 r0 *1 28.2,5.98
X$121 161 162 163 7 164 10 257 258 cell_2rw
* cell instance $122 r0 *1 29.375,5.98
X$122 165 166 167 7 168 10 257 258 cell_2rw
* cell instance $123 r0 *1 30.55,5.98
X$123 169 170 171 7 172 10 257 258 cell_2rw
* cell instance $124 r0 *1 31.725,5.98
X$124 173 174 175 7 176 10 257 258 cell_2rw
* cell instance $125 r0 *1 32.9,5.98
X$125 177 178 179 7 180 10 257 258 cell_2rw
* cell instance $126 r0 *1 34.075,5.98
X$126 181 182 183 7 184 10 257 258 cell_2rw
* cell instance $127 r0 *1 35.25,5.98
X$127 185 186 187 7 188 10 257 258 cell_2rw
* cell instance $128 r0 *1 36.425,5.98
X$128 189 190 191 7 192 10 257 258 cell_2rw
* cell instance $129 m0 *1 1.175,8.97
X$129 65 66 67 9 68 8 257 258 cell_2rw
* cell instance $130 m0 *1 0,8.97
X$130 61 62 63 9 64 8 257 258 cell_2rw
* cell instance $131 m0 *1 2.35,8.97
X$131 69 70 71 9 72 8 257 258 cell_2rw
* cell instance $132 m0 *1 3.525,8.97
X$132 73 74 75 9 76 8 257 258 cell_2rw
* cell instance $133 m0 *1 4.7,8.97
X$133 77 78 79 9 80 8 257 258 cell_2rw
* cell instance $134 m0 *1 5.875,8.97
X$134 81 82 83 9 84 8 257 258 cell_2rw
* cell instance $135 m0 *1 7.05,8.97
X$135 85 86 87 9 88 8 257 258 cell_2rw
* cell instance $136 m0 *1 8.225,8.97
X$136 89 90 91 9 92 8 257 258 cell_2rw
* cell instance $137 m0 *1 9.4,8.97
X$137 93 94 95 9 96 8 257 258 cell_2rw
* cell instance $138 m0 *1 10.575,8.97
X$138 97 98 99 9 100 8 257 258 cell_2rw
* cell instance $139 m0 *1 11.75,8.97
X$139 101 102 103 9 104 8 257 258 cell_2rw
* cell instance $140 m0 *1 12.925,8.97
X$140 105 106 107 9 108 8 257 258 cell_2rw
* cell instance $141 m0 *1 14.1,8.97
X$141 109 110 111 9 112 8 257 258 cell_2rw
* cell instance $142 m0 *1 15.275,8.97
X$142 113 114 115 9 116 8 257 258 cell_2rw
* cell instance $143 m0 *1 16.45,8.97
X$143 117 118 119 9 120 8 257 258 cell_2rw
* cell instance $144 m0 *1 17.625,8.97
X$144 121 122 123 9 124 8 257 258 cell_2rw
* cell instance $145 m0 *1 18.8,8.97
X$145 129 130 131 9 132 8 257 258 cell_2rw
* cell instance $146 m0 *1 19.975,8.97
X$146 133 134 135 9 136 8 257 258 cell_2rw
* cell instance $147 m0 *1 21.15,8.97
X$147 137 138 139 9 140 8 257 258 cell_2rw
* cell instance $148 m0 *1 22.325,8.97
X$148 141 142 143 9 144 8 257 258 cell_2rw
* cell instance $149 m0 *1 23.5,8.97
X$149 145 146 147 9 148 8 257 258 cell_2rw
* cell instance $150 m0 *1 24.675,8.97
X$150 149 150 151 9 152 8 257 258 cell_2rw
* cell instance $151 m0 *1 25.85,8.97
X$151 153 154 155 9 156 8 257 258 cell_2rw
* cell instance $152 m0 *1 27.025,8.97
X$152 157 158 159 9 160 8 257 258 cell_2rw
* cell instance $153 m0 *1 28.2,8.97
X$153 161 162 163 9 164 8 257 258 cell_2rw
* cell instance $154 m0 *1 29.375,8.97
X$154 165 166 167 9 168 8 257 258 cell_2rw
* cell instance $155 m0 *1 30.55,8.97
X$155 169 170 171 9 172 8 257 258 cell_2rw
* cell instance $156 m0 *1 31.725,8.97
X$156 173 174 175 9 176 8 257 258 cell_2rw
* cell instance $157 m0 *1 32.9,8.97
X$157 177 178 179 9 180 8 257 258 cell_2rw
* cell instance $158 m0 *1 34.075,8.97
X$158 181 182 183 9 184 8 257 258 cell_2rw
* cell instance $159 m0 *1 35.25,8.97
X$159 185 186 187 9 188 8 257 258 cell_2rw
* cell instance $160 m0 *1 36.425,8.97
X$160 189 190 191 9 192 8 257 258 cell_2rw
* cell instance $161 m0 *1 1.175,5.98
X$161 65 66 67 11 68 12 257 258 cell_2rw
* cell instance $162 m0 *1 0,5.98
X$162 61 62 63 11 64 12 257 258 cell_2rw
* cell instance $163 m0 *1 2.35,5.98
X$163 69 70 71 11 72 12 257 258 cell_2rw
* cell instance $164 m0 *1 3.525,5.98
X$164 73 74 75 11 76 12 257 258 cell_2rw
* cell instance $165 m0 *1 4.7,5.98
X$165 77 78 79 11 80 12 257 258 cell_2rw
* cell instance $166 m0 *1 5.875,5.98
X$166 81 82 83 11 84 12 257 258 cell_2rw
* cell instance $167 m0 *1 7.05,5.98
X$167 85 86 87 11 88 12 257 258 cell_2rw
* cell instance $168 m0 *1 8.225,5.98
X$168 89 90 91 11 92 12 257 258 cell_2rw
* cell instance $169 m0 *1 9.4,5.98
X$169 93 94 95 11 96 12 257 258 cell_2rw
* cell instance $170 m0 *1 10.575,5.98
X$170 97 98 99 11 100 12 257 258 cell_2rw
* cell instance $171 m0 *1 11.75,5.98
X$171 101 102 103 11 104 12 257 258 cell_2rw
* cell instance $172 m0 *1 12.925,5.98
X$172 105 106 107 11 108 12 257 258 cell_2rw
* cell instance $173 m0 *1 14.1,5.98
X$173 109 110 111 11 112 12 257 258 cell_2rw
* cell instance $174 m0 *1 15.275,5.98
X$174 113 114 115 11 116 12 257 258 cell_2rw
* cell instance $175 m0 *1 16.45,5.98
X$175 117 118 119 11 120 12 257 258 cell_2rw
* cell instance $176 m0 *1 17.625,5.98
X$176 121 122 123 11 124 12 257 258 cell_2rw
* cell instance $177 m0 *1 18.8,5.98
X$177 129 130 131 11 132 12 257 258 cell_2rw
* cell instance $178 m0 *1 19.975,5.98
X$178 133 134 135 11 136 12 257 258 cell_2rw
* cell instance $179 m0 *1 21.15,5.98
X$179 137 138 139 11 140 12 257 258 cell_2rw
* cell instance $180 m0 *1 22.325,5.98
X$180 141 142 143 11 144 12 257 258 cell_2rw
* cell instance $181 m0 *1 23.5,5.98
X$181 145 146 147 11 148 12 257 258 cell_2rw
* cell instance $182 m0 *1 24.675,5.98
X$182 149 150 151 11 152 12 257 258 cell_2rw
* cell instance $183 m0 *1 25.85,5.98
X$183 153 154 155 11 156 12 257 258 cell_2rw
* cell instance $184 m0 *1 27.025,5.98
X$184 157 158 159 11 160 12 257 258 cell_2rw
* cell instance $185 m0 *1 28.2,5.98
X$185 161 162 163 11 164 12 257 258 cell_2rw
* cell instance $186 m0 *1 29.375,5.98
X$186 165 166 167 11 168 12 257 258 cell_2rw
* cell instance $187 m0 *1 30.55,5.98
X$187 169 170 171 11 172 12 257 258 cell_2rw
* cell instance $188 m0 *1 31.725,5.98
X$188 173 174 175 11 176 12 257 258 cell_2rw
* cell instance $189 m0 *1 32.9,5.98
X$189 177 178 179 11 180 12 257 258 cell_2rw
* cell instance $190 m0 *1 34.075,5.98
X$190 181 182 183 11 184 12 257 258 cell_2rw
* cell instance $191 m0 *1 35.25,5.98
X$191 185 186 187 11 188 12 257 258 cell_2rw
* cell instance $192 m0 *1 36.425,5.98
X$192 189 190 191 11 192 12 257 258 cell_2rw
* cell instance $193 m0 *1 1.175,11.96
X$193 65 66 67 13 68 14 257 258 cell_2rw
* cell instance $194 m0 *1 0,11.96
X$194 61 62 63 13 64 14 257 258 cell_2rw
* cell instance $195 m0 *1 2.35,11.96
X$195 69 70 71 13 72 14 257 258 cell_2rw
* cell instance $196 m0 *1 3.525,11.96
X$196 73 74 75 13 76 14 257 258 cell_2rw
* cell instance $197 m0 *1 4.7,11.96
X$197 77 78 79 13 80 14 257 258 cell_2rw
* cell instance $198 m0 *1 5.875,11.96
X$198 81 82 83 13 84 14 257 258 cell_2rw
* cell instance $199 m0 *1 7.05,11.96
X$199 85 86 87 13 88 14 257 258 cell_2rw
* cell instance $200 m0 *1 8.225,11.96
X$200 89 90 91 13 92 14 257 258 cell_2rw
* cell instance $201 m0 *1 9.4,11.96
X$201 93 94 95 13 96 14 257 258 cell_2rw
* cell instance $202 m0 *1 10.575,11.96
X$202 97 98 99 13 100 14 257 258 cell_2rw
* cell instance $203 m0 *1 11.75,11.96
X$203 101 102 103 13 104 14 257 258 cell_2rw
* cell instance $204 m0 *1 12.925,11.96
X$204 105 106 107 13 108 14 257 258 cell_2rw
* cell instance $205 m0 *1 14.1,11.96
X$205 109 110 111 13 112 14 257 258 cell_2rw
* cell instance $206 m0 *1 15.275,11.96
X$206 113 114 115 13 116 14 257 258 cell_2rw
* cell instance $207 m0 *1 16.45,11.96
X$207 117 118 119 13 120 14 257 258 cell_2rw
* cell instance $208 m0 *1 17.625,11.96
X$208 121 122 123 13 124 14 257 258 cell_2rw
* cell instance $209 m0 *1 18.8,11.96
X$209 129 130 131 13 132 14 257 258 cell_2rw
* cell instance $210 m0 *1 19.975,11.96
X$210 133 134 135 13 136 14 257 258 cell_2rw
* cell instance $211 m0 *1 21.15,11.96
X$211 137 138 139 13 140 14 257 258 cell_2rw
* cell instance $212 m0 *1 22.325,11.96
X$212 141 142 143 13 144 14 257 258 cell_2rw
* cell instance $213 m0 *1 23.5,11.96
X$213 145 146 147 13 148 14 257 258 cell_2rw
* cell instance $214 m0 *1 24.675,11.96
X$214 149 150 151 13 152 14 257 258 cell_2rw
* cell instance $215 m0 *1 25.85,11.96
X$215 153 154 155 13 156 14 257 258 cell_2rw
* cell instance $216 m0 *1 27.025,11.96
X$216 157 158 159 13 160 14 257 258 cell_2rw
* cell instance $217 m0 *1 28.2,11.96
X$217 161 162 163 13 164 14 257 258 cell_2rw
* cell instance $218 m0 *1 29.375,11.96
X$218 165 166 167 13 168 14 257 258 cell_2rw
* cell instance $219 m0 *1 30.55,11.96
X$219 169 170 171 13 172 14 257 258 cell_2rw
* cell instance $220 m0 *1 31.725,11.96
X$220 173 174 175 13 176 14 257 258 cell_2rw
* cell instance $221 m0 *1 32.9,11.96
X$221 177 178 179 13 180 14 257 258 cell_2rw
* cell instance $222 m0 *1 34.075,11.96
X$222 181 182 183 13 184 14 257 258 cell_2rw
* cell instance $223 m0 *1 35.25,11.96
X$223 185 186 187 13 188 14 257 258 cell_2rw
* cell instance $224 m0 *1 36.425,11.96
X$224 189 190 191 13 192 14 257 258 cell_2rw
* cell instance $225 r0 *1 1.175,11.96
X$225 65 66 67 16 68 15 257 258 cell_2rw
* cell instance $226 r0 *1 0,11.96
X$226 61 62 63 16 64 15 257 258 cell_2rw
* cell instance $227 r0 *1 2.35,11.96
X$227 69 70 71 16 72 15 257 258 cell_2rw
* cell instance $228 r0 *1 3.525,11.96
X$228 73 74 75 16 76 15 257 258 cell_2rw
* cell instance $229 r0 *1 4.7,11.96
X$229 77 78 79 16 80 15 257 258 cell_2rw
* cell instance $230 r0 *1 5.875,11.96
X$230 81 82 83 16 84 15 257 258 cell_2rw
* cell instance $231 r0 *1 7.05,11.96
X$231 85 86 87 16 88 15 257 258 cell_2rw
* cell instance $232 r0 *1 8.225,11.96
X$232 89 90 91 16 92 15 257 258 cell_2rw
* cell instance $233 r0 *1 9.4,11.96
X$233 93 94 95 16 96 15 257 258 cell_2rw
* cell instance $234 r0 *1 10.575,11.96
X$234 97 98 99 16 100 15 257 258 cell_2rw
* cell instance $235 r0 *1 11.75,11.96
X$235 101 102 103 16 104 15 257 258 cell_2rw
* cell instance $236 r0 *1 12.925,11.96
X$236 105 106 107 16 108 15 257 258 cell_2rw
* cell instance $237 r0 *1 14.1,11.96
X$237 109 110 111 16 112 15 257 258 cell_2rw
* cell instance $238 r0 *1 15.275,11.96
X$238 113 114 115 16 116 15 257 258 cell_2rw
* cell instance $239 r0 *1 16.45,11.96
X$239 117 118 119 16 120 15 257 258 cell_2rw
* cell instance $240 r0 *1 17.625,11.96
X$240 121 122 123 16 124 15 257 258 cell_2rw
* cell instance $241 r0 *1 18.8,11.96
X$241 129 130 131 16 132 15 257 258 cell_2rw
* cell instance $242 r0 *1 19.975,11.96
X$242 133 134 135 16 136 15 257 258 cell_2rw
* cell instance $243 r0 *1 21.15,11.96
X$243 137 138 139 16 140 15 257 258 cell_2rw
* cell instance $244 r0 *1 22.325,11.96
X$244 141 142 143 16 144 15 257 258 cell_2rw
* cell instance $245 r0 *1 23.5,11.96
X$245 145 146 147 16 148 15 257 258 cell_2rw
* cell instance $246 r0 *1 24.675,11.96
X$246 149 150 151 16 152 15 257 258 cell_2rw
* cell instance $247 r0 *1 25.85,11.96
X$247 153 154 155 16 156 15 257 258 cell_2rw
* cell instance $248 r0 *1 27.025,11.96
X$248 157 158 159 16 160 15 257 258 cell_2rw
* cell instance $249 r0 *1 28.2,11.96
X$249 161 162 163 16 164 15 257 258 cell_2rw
* cell instance $250 r0 *1 29.375,11.96
X$250 165 166 167 16 168 15 257 258 cell_2rw
* cell instance $251 r0 *1 30.55,11.96
X$251 169 170 171 16 172 15 257 258 cell_2rw
* cell instance $252 r0 *1 31.725,11.96
X$252 173 174 175 16 176 15 257 258 cell_2rw
* cell instance $253 r0 *1 32.9,11.96
X$253 177 178 179 16 180 15 257 258 cell_2rw
* cell instance $254 r0 *1 34.075,11.96
X$254 181 182 183 16 184 15 257 258 cell_2rw
* cell instance $255 r0 *1 35.25,11.96
X$255 185 186 187 16 188 15 257 258 cell_2rw
* cell instance $256 r0 *1 36.425,11.96
X$256 189 190 191 16 192 15 257 258 cell_2rw
* cell instance $257 r0 *1 1.175,8.97
X$257 65 66 67 17 68 18 257 258 cell_2rw
* cell instance $258 r0 *1 0,8.97
X$258 61 62 63 17 64 18 257 258 cell_2rw
* cell instance $259 r0 *1 2.35,8.97
X$259 69 70 71 17 72 18 257 258 cell_2rw
* cell instance $260 r0 *1 3.525,8.97
X$260 73 74 75 17 76 18 257 258 cell_2rw
* cell instance $261 r0 *1 4.7,8.97
X$261 77 78 79 17 80 18 257 258 cell_2rw
* cell instance $262 r0 *1 5.875,8.97
X$262 81 82 83 17 84 18 257 258 cell_2rw
* cell instance $263 r0 *1 7.05,8.97
X$263 85 86 87 17 88 18 257 258 cell_2rw
* cell instance $264 r0 *1 8.225,8.97
X$264 89 90 91 17 92 18 257 258 cell_2rw
* cell instance $265 r0 *1 9.4,8.97
X$265 93 94 95 17 96 18 257 258 cell_2rw
* cell instance $266 r0 *1 10.575,8.97
X$266 97 98 99 17 100 18 257 258 cell_2rw
* cell instance $267 r0 *1 11.75,8.97
X$267 101 102 103 17 104 18 257 258 cell_2rw
* cell instance $268 r0 *1 12.925,8.97
X$268 105 106 107 17 108 18 257 258 cell_2rw
* cell instance $269 r0 *1 14.1,8.97
X$269 109 110 111 17 112 18 257 258 cell_2rw
* cell instance $270 r0 *1 15.275,8.97
X$270 113 114 115 17 116 18 257 258 cell_2rw
* cell instance $271 r0 *1 16.45,8.97
X$271 117 118 119 17 120 18 257 258 cell_2rw
* cell instance $272 r0 *1 17.625,8.97
X$272 121 122 123 17 124 18 257 258 cell_2rw
* cell instance $273 r0 *1 18.8,8.97
X$273 129 130 131 17 132 18 257 258 cell_2rw
* cell instance $274 r0 *1 19.975,8.97
X$274 133 134 135 17 136 18 257 258 cell_2rw
* cell instance $275 r0 *1 21.15,8.97
X$275 137 138 139 17 140 18 257 258 cell_2rw
* cell instance $276 r0 *1 22.325,8.97
X$276 141 142 143 17 144 18 257 258 cell_2rw
* cell instance $277 r0 *1 23.5,8.97
X$277 145 146 147 17 148 18 257 258 cell_2rw
* cell instance $278 r0 *1 24.675,8.97
X$278 149 150 151 17 152 18 257 258 cell_2rw
* cell instance $279 r0 *1 25.85,8.97
X$279 153 154 155 17 156 18 257 258 cell_2rw
* cell instance $280 r0 *1 27.025,8.97
X$280 157 158 159 17 160 18 257 258 cell_2rw
* cell instance $281 r0 *1 28.2,8.97
X$281 161 162 163 17 164 18 257 258 cell_2rw
* cell instance $282 r0 *1 29.375,8.97
X$282 165 166 167 17 168 18 257 258 cell_2rw
* cell instance $283 r0 *1 30.55,8.97
X$283 169 170 171 17 172 18 257 258 cell_2rw
* cell instance $284 r0 *1 31.725,8.97
X$284 173 174 175 17 176 18 257 258 cell_2rw
* cell instance $285 r0 *1 32.9,8.97
X$285 177 178 179 17 180 18 257 258 cell_2rw
* cell instance $286 r0 *1 34.075,8.97
X$286 181 182 183 17 184 18 257 258 cell_2rw
* cell instance $287 r0 *1 35.25,8.97
X$287 185 186 187 17 188 18 257 258 cell_2rw
* cell instance $288 r0 *1 36.425,8.97
X$288 189 190 191 17 192 18 257 258 cell_2rw
* cell instance $289 r0 *1 1.175,14.95
X$289 65 66 67 20 68 19 257 258 cell_2rw
* cell instance $290 r0 *1 0,14.95
X$290 61 62 63 20 64 19 257 258 cell_2rw
* cell instance $291 r0 *1 2.35,14.95
X$291 69 70 71 20 72 19 257 258 cell_2rw
* cell instance $292 r0 *1 3.525,14.95
X$292 73 74 75 20 76 19 257 258 cell_2rw
* cell instance $293 r0 *1 4.7,14.95
X$293 77 78 79 20 80 19 257 258 cell_2rw
* cell instance $294 r0 *1 5.875,14.95
X$294 81 82 83 20 84 19 257 258 cell_2rw
* cell instance $295 r0 *1 7.05,14.95
X$295 85 86 87 20 88 19 257 258 cell_2rw
* cell instance $296 r0 *1 8.225,14.95
X$296 89 90 91 20 92 19 257 258 cell_2rw
* cell instance $297 r0 *1 9.4,14.95
X$297 93 94 95 20 96 19 257 258 cell_2rw
* cell instance $298 r0 *1 10.575,14.95
X$298 97 98 99 20 100 19 257 258 cell_2rw
* cell instance $299 r0 *1 11.75,14.95
X$299 101 102 103 20 104 19 257 258 cell_2rw
* cell instance $300 r0 *1 12.925,14.95
X$300 105 106 107 20 108 19 257 258 cell_2rw
* cell instance $301 r0 *1 14.1,14.95
X$301 109 110 111 20 112 19 257 258 cell_2rw
* cell instance $302 r0 *1 15.275,14.95
X$302 113 114 115 20 116 19 257 258 cell_2rw
* cell instance $303 r0 *1 16.45,14.95
X$303 117 118 119 20 120 19 257 258 cell_2rw
* cell instance $304 r0 *1 17.625,14.95
X$304 121 122 123 20 124 19 257 258 cell_2rw
* cell instance $305 r0 *1 18.8,14.95
X$305 129 130 131 20 132 19 257 258 cell_2rw
* cell instance $306 r0 *1 19.975,14.95
X$306 133 134 135 20 136 19 257 258 cell_2rw
* cell instance $307 r0 *1 21.15,14.95
X$307 137 138 139 20 140 19 257 258 cell_2rw
* cell instance $308 r0 *1 22.325,14.95
X$308 141 142 143 20 144 19 257 258 cell_2rw
* cell instance $309 r0 *1 23.5,14.95
X$309 145 146 147 20 148 19 257 258 cell_2rw
* cell instance $310 r0 *1 24.675,14.95
X$310 149 150 151 20 152 19 257 258 cell_2rw
* cell instance $311 r0 *1 25.85,14.95
X$311 153 154 155 20 156 19 257 258 cell_2rw
* cell instance $312 r0 *1 27.025,14.95
X$312 157 158 159 20 160 19 257 258 cell_2rw
* cell instance $313 r0 *1 28.2,14.95
X$313 161 162 163 20 164 19 257 258 cell_2rw
* cell instance $314 r0 *1 29.375,14.95
X$314 165 166 167 20 168 19 257 258 cell_2rw
* cell instance $315 r0 *1 30.55,14.95
X$315 169 170 171 20 172 19 257 258 cell_2rw
* cell instance $316 r0 *1 31.725,14.95
X$316 173 174 175 20 176 19 257 258 cell_2rw
* cell instance $317 r0 *1 32.9,14.95
X$317 177 178 179 20 180 19 257 258 cell_2rw
* cell instance $318 r0 *1 34.075,14.95
X$318 181 182 183 20 184 19 257 258 cell_2rw
* cell instance $319 r0 *1 35.25,14.95
X$319 185 186 187 20 188 19 257 258 cell_2rw
* cell instance $320 r0 *1 36.425,14.95
X$320 189 190 191 20 192 19 257 258 cell_2rw
* cell instance $321 m0 *1 1.175,17.94
X$321 65 66 67 21 68 22 257 258 cell_2rw
* cell instance $322 m0 *1 0,17.94
X$322 61 62 63 21 64 22 257 258 cell_2rw
* cell instance $323 m0 *1 2.35,17.94
X$323 69 70 71 21 72 22 257 258 cell_2rw
* cell instance $324 m0 *1 3.525,17.94
X$324 73 74 75 21 76 22 257 258 cell_2rw
* cell instance $325 m0 *1 4.7,17.94
X$325 77 78 79 21 80 22 257 258 cell_2rw
* cell instance $326 m0 *1 5.875,17.94
X$326 81 82 83 21 84 22 257 258 cell_2rw
* cell instance $327 m0 *1 7.05,17.94
X$327 85 86 87 21 88 22 257 258 cell_2rw
* cell instance $328 m0 *1 8.225,17.94
X$328 89 90 91 21 92 22 257 258 cell_2rw
* cell instance $329 m0 *1 9.4,17.94
X$329 93 94 95 21 96 22 257 258 cell_2rw
* cell instance $330 m0 *1 10.575,17.94
X$330 97 98 99 21 100 22 257 258 cell_2rw
* cell instance $331 m0 *1 11.75,17.94
X$331 101 102 103 21 104 22 257 258 cell_2rw
* cell instance $332 m0 *1 12.925,17.94
X$332 105 106 107 21 108 22 257 258 cell_2rw
* cell instance $333 m0 *1 14.1,17.94
X$333 109 110 111 21 112 22 257 258 cell_2rw
* cell instance $334 m0 *1 15.275,17.94
X$334 113 114 115 21 116 22 257 258 cell_2rw
* cell instance $335 m0 *1 16.45,17.94
X$335 117 118 119 21 120 22 257 258 cell_2rw
* cell instance $336 m0 *1 17.625,17.94
X$336 121 122 123 21 124 22 257 258 cell_2rw
* cell instance $337 m0 *1 18.8,17.94
X$337 129 130 131 21 132 22 257 258 cell_2rw
* cell instance $338 m0 *1 19.975,17.94
X$338 133 134 135 21 136 22 257 258 cell_2rw
* cell instance $339 m0 *1 21.15,17.94
X$339 137 138 139 21 140 22 257 258 cell_2rw
* cell instance $340 m0 *1 22.325,17.94
X$340 141 142 143 21 144 22 257 258 cell_2rw
* cell instance $341 m0 *1 23.5,17.94
X$341 145 146 147 21 148 22 257 258 cell_2rw
* cell instance $342 m0 *1 24.675,17.94
X$342 149 150 151 21 152 22 257 258 cell_2rw
* cell instance $343 m0 *1 25.85,17.94
X$343 153 154 155 21 156 22 257 258 cell_2rw
* cell instance $344 m0 *1 27.025,17.94
X$344 157 158 159 21 160 22 257 258 cell_2rw
* cell instance $345 m0 *1 28.2,17.94
X$345 161 162 163 21 164 22 257 258 cell_2rw
* cell instance $346 m0 *1 29.375,17.94
X$346 165 166 167 21 168 22 257 258 cell_2rw
* cell instance $347 m0 *1 30.55,17.94
X$347 169 170 171 21 172 22 257 258 cell_2rw
* cell instance $348 m0 *1 31.725,17.94
X$348 173 174 175 21 176 22 257 258 cell_2rw
* cell instance $349 m0 *1 32.9,17.94
X$349 177 178 179 21 180 22 257 258 cell_2rw
* cell instance $350 m0 *1 34.075,17.94
X$350 181 182 183 21 184 22 257 258 cell_2rw
* cell instance $351 m0 *1 35.25,17.94
X$351 185 186 187 21 188 22 257 258 cell_2rw
* cell instance $352 m0 *1 36.425,17.94
X$352 189 190 191 21 192 22 257 258 cell_2rw
* cell instance $353 m0 *1 1.175,14.95
X$353 65 66 67 24 68 23 257 258 cell_2rw
* cell instance $354 m0 *1 0,14.95
X$354 61 62 63 24 64 23 257 258 cell_2rw
* cell instance $355 m0 *1 2.35,14.95
X$355 69 70 71 24 72 23 257 258 cell_2rw
* cell instance $356 m0 *1 3.525,14.95
X$356 73 74 75 24 76 23 257 258 cell_2rw
* cell instance $357 m0 *1 4.7,14.95
X$357 77 78 79 24 80 23 257 258 cell_2rw
* cell instance $358 m0 *1 5.875,14.95
X$358 81 82 83 24 84 23 257 258 cell_2rw
* cell instance $359 m0 *1 7.05,14.95
X$359 85 86 87 24 88 23 257 258 cell_2rw
* cell instance $360 m0 *1 8.225,14.95
X$360 89 90 91 24 92 23 257 258 cell_2rw
* cell instance $361 m0 *1 9.4,14.95
X$361 93 94 95 24 96 23 257 258 cell_2rw
* cell instance $362 m0 *1 10.575,14.95
X$362 97 98 99 24 100 23 257 258 cell_2rw
* cell instance $363 m0 *1 11.75,14.95
X$363 101 102 103 24 104 23 257 258 cell_2rw
* cell instance $364 m0 *1 12.925,14.95
X$364 105 106 107 24 108 23 257 258 cell_2rw
* cell instance $365 m0 *1 14.1,14.95
X$365 109 110 111 24 112 23 257 258 cell_2rw
* cell instance $366 m0 *1 15.275,14.95
X$366 113 114 115 24 116 23 257 258 cell_2rw
* cell instance $367 m0 *1 16.45,14.95
X$367 117 118 119 24 120 23 257 258 cell_2rw
* cell instance $368 m0 *1 17.625,14.95
X$368 121 122 123 24 124 23 257 258 cell_2rw
* cell instance $369 m0 *1 18.8,14.95
X$369 129 130 131 24 132 23 257 258 cell_2rw
* cell instance $370 m0 *1 19.975,14.95
X$370 133 134 135 24 136 23 257 258 cell_2rw
* cell instance $371 m0 *1 21.15,14.95
X$371 137 138 139 24 140 23 257 258 cell_2rw
* cell instance $372 m0 *1 22.325,14.95
X$372 141 142 143 24 144 23 257 258 cell_2rw
* cell instance $373 m0 *1 23.5,14.95
X$373 145 146 147 24 148 23 257 258 cell_2rw
* cell instance $374 m0 *1 24.675,14.95
X$374 149 150 151 24 152 23 257 258 cell_2rw
* cell instance $375 m0 *1 25.85,14.95
X$375 153 154 155 24 156 23 257 258 cell_2rw
* cell instance $376 m0 *1 27.025,14.95
X$376 157 158 159 24 160 23 257 258 cell_2rw
* cell instance $377 m0 *1 28.2,14.95
X$377 161 162 163 24 164 23 257 258 cell_2rw
* cell instance $378 m0 *1 29.375,14.95
X$378 165 166 167 24 168 23 257 258 cell_2rw
* cell instance $379 m0 *1 30.55,14.95
X$379 169 170 171 24 172 23 257 258 cell_2rw
* cell instance $380 m0 *1 31.725,14.95
X$380 173 174 175 24 176 23 257 258 cell_2rw
* cell instance $381 m0 *1 32.9,14.95
X$381 177 178 179 24 180 23 257 258 cell_2rw
* cell instance $382 m0 *1 34.075,14.95
X$382 181 182 183 24 184 23 257 258 cell_2rw
* cell instance $383 m0 *1 35.25,14.95
X$383 185 186 187 24 188 23 257 258 cell_2rw
* cell instance $384 m0 *1 36.425,14.95
X$384 189 190 191 24 192 23 257 258 cell_2rw
* cell instance $385 r0 *1 1.175,20.93
X$385 65 66 67 28 68 25 257 258 cell_2rw
* cell instance $386 r0 *1 0,20.93
X$386 61 62 63 28 64 25 257 258 cell_2rw
* cell instance $387 r0 *1 2.35,20.93
X$387 69 70 71 28 72 25 257 258 cell_2rw
* cell instance $388 r0 *1 3.525,20.93
X$388 73 74 75 28 76 25 257 258 cell_2rw
* cell instance $389 r0 *1 4.7,20.93
X$389 77 78 79 28 80 25 257 258 cell_2rw
* cell instance $390 r0 *1 5.875,20.93
X$390 81 82 83 28 84 25 257 258 cell_2rw
* cell instance $391 r0 *1 7.05,20.93
X$391 85 86 87 28 88 25 257 258 cell_2rw
* cell instance $392 r0 *1 8.225,20.93
X$392 89 90 91 28 92 25 257 258 cell_2rw
* cell instance $393 r0 *1 9.4,20.93
X$393 93 94 95 28 96 25 257 258 cell_2rw
* cell instance $394 r0 *1 10.575,20.93
X$394 97 98 99 28 100 25 257 258 cell_2rw
* cell instance $395 r0 *1 11.75,20.93
X$395 101 102 103 28 104 25 257 258 cell_2rw
* cell instance $396 r0 *1 12.925,20.93
X$396 105 106 107 28 108 25 257 258 cell_2rw
* cell instance $397 r0 *1 14.1,20.93
X$397 109 110 111 28 112 25 257 258 cell_2rw
* cell instance $398 r0 *1 15.275,20.93
X$398 113 114 115 28 116 25 257 258 cell_2rw
* cell instance $399 r0 *1 16.45,20.93
X$399 117 118 119 28 120 25 257 258 cell_2rw
* cell instance $400 r0 *1 17.625,20.93
X$400 121 122 123 28 124 25 257 258 cell_2rw
* cell instance $401 r0 *1 18.8,20.93
X$401 129 130 131 28 132 25 257 258 cell_2rw
* cell instance $402 r0 *1 19.975,20.93
X$402 133 134 135 28 136 25 257 258 cell_2rw
* cell instance $403 r0 *1 21.15,20.93
X$403 137 138 139 28 140 25 257 258 cell_2rw
* cell instance $404 r0 *1 22.325,20.93
X$404 141 142 143 28 144 25 257 258 cell_2rw
* cell instance $405 r0 *1 23.5,20.93
X$405 145 146 147 28 148 25 257 258 cell_2rw
* cell instance $406 r0 *1 24.675,20.93
X$406 149 150 151 28 152 25 257 258 cell_2rw
* cell instance $407 r0 *1 25.85,20.93
X$407 153 154 155 28 156 25 257 258 cell_2rw
* cell instance $408 r0 *1 27.025,20.93
X$408 157 158 159 28 160 25 257 258 cell_2rw
* cell instance $409 r0 *1 28.2,20.93
X$409 161 162 163 28 164 25 257 258 cell_2rw
* cell instance $410 r0 *1 29.375,20.93
X$410 165 166 167 28 168 25 257 258 cell_2rw
* cell instance $411 r0 *1 30.55,20.93
X$411 169 170 171 28 172 25 257 258 cell_2rw
* cell instance $412 r0 *1 31.725,20.93
X$412 173 174 175 28 176 25 257 258 cell_2rw
* cell instance $413 r0 *1 32.9,20.93
X$413 177 178 179 28 180 25 257 258 cell_2rw
* cell instance $414 r0 *1 34.075,20.93
X$414 181 182 183 28 184 25 257 258 cell_2rw
* cell instance $415 r0 *1 35.25,20.93
X$415 185 186 187 28 188 25 257 258 cell_2rw
* cell instance $416 r0 *1 36.425,20.93
X$416 189 190 191 28 192 25 257 258 cell_2rw
* cell instance $417 m0 *1 1.175,20.93
X$417 65 66 67 26 68 29 257 258 cell_2rw
* cell instance $418 m0 *1 0,20.93
X$418 61 62 63 26 64 29 257 258 cell_2rw
* cell instance $419 m0 *1 2.35,20.93
X$419 69 70 71 26 72 29 257 258 cell_2rw
* cell instance $420 m0 *1 3.525,20.93
X$420 73 74 75 26 76 29 257 258 cell_2rw
* cell instance $421 m0 *1 4.7,20.93
X$421 77 78 79 26 80 29 257 258 cell_2rw
* cell instance $422 m0 *1 5.875,20.93
X$422 81 82 83 26 84 29 257 258 cell_2rw
* cell instance $423 m0 *1 7.05,20.93
X$423 85 86 87 26 88 29 257 258 cell_2rw
* cell instance $424 m0 *1 8.225,20.93
X$424 89 90 91 26 92 29 257 258 cell_2rw
* cell instance $425 m0 *1 9.4,20.93
X$425 93 94 95 26 96 29 257 258 cell_2rw
* cell instance $426 m0 *1 10.575,20.93
X$426 97 98 99 26 100 29 257 258 cell_2rw
* cell instance $427 m0 *1 11.75,20.93
X$427 101 102 103 26 104 29 257 258 cell_2rw
* cell instance $428 m0 *1 12.925,20.93
X$428 105 106 107 26 108 29 257 258 cell_2rw
* cell instance $429 m0 *1 14.1,20.93
X$429 109 110 111 26 112 29 257 258 cell_2rw
* cell instance $430 m0 *1 15.275,20.93
X$430 113 114 115 26 116 29 257 258 cell_2rw
* cell instance $431 m0 *1 16.45,20.93
X$431 117 118 119 26 120 29 257 258 cell_2rw
* cell instance $432 m0 *1 17.625,20.93
X$432 121 122 123 26 124 29 257 258 cell_2rw
* cell instance $433 m0 *1 18.8,20.93
X$433 129 130 131 26 132 29 257 258 cell_2rw
* cell instance $434 m0 *1 19.975,20.93
X$434 133 134 135 26 136 29 257 258 cell_2rw
* cell instance $435 m0 *1 21.15,20.93
X$435 137 138 139 26 140 29 257 258 cell_2rw
* cell instance $436 m0 *1 22.325,20.93
X$436 141 142 143 26 144 29 257 258 cell_2rw
* cell instance $437 m0 *1 23.5,20.93
X$437 145 146 147 26 148 29 257 258 cell_2rw
* cell instance $438 m0 *1 24.675,20.93
X$438 149 150 151 26 152 29 257 258 cell_2rw
* cell instance $439 m0 *1 25.85,20.93
X$439 153 154 155 26 156 29 257 258 cell_2rw
* cell instance $440 m0 *1 27.025,20.93
X$440 157 158 159 26 160 29 257 258 cell_2rw
* cell instance $441 m0 *1 28.2,20.93
X$441 161 162 163 26 164 29 257 258 cell_2rw
* cell instance $442 m0 *1 29.375,20.93
X$442 165 166 167 26 168 29 257 258 cell_2rw
* cell instance $443 m0 *1 30.55,20.93
X$443 169 170 171 26 172 29 257 258 cell_2rw
* cell instance $444 m0 *1 31.725,20.93
X$444 173 174 175 26 176 29 257 258 cell_2rw
* cell instance $445 m0 *1 32.9,20.93
X$445 177 178 179 26 180 29 257 258 cell_2rw
* cell instance $446 m0 *1 34.075,20.93
X$446 181 182 183 26 184 29 257 258 cell_2rw
* cell instance $447 m0 *1 35.25,20.93
X$447 185 186 187 26 188 29 257 258 cell_2rw
* cell instance $448 m0 *1 36.425,20.93
X$448 189 190 191 26 192 29 257 258 cell_2rw
* cell instance $449 r0 *1 1.175,17.94
X$449 65 66 67 27 68 30 257 258 cell_2rw
* cell instance $450 r0 *1 0,17.94
X$450 61 62 63 27 64 30 257 258 cell_2rw
* cell instance $451 r0 *1 2.35,17.94
X$451 69 70 71 27 72 30 257 258 cell_2rw
* cell instance $452 r0 *1 3.525,17.94
X$452 73 74 75 27 76 30 257 258 cell_2rw
* cell instance $453 r0 *1 4.7,17.94
X$453 77 78 79 27 80 30 257 258 cell_2rw
* cell instance $454 r0 *1 5.875,17.94
X$454 81 82 83 27 84 30 257 258 cell_2rw
* cell instance $455 r0 *1 7.05,17.94
X$455 85 86 87 27 88 30 257 258 cell_2rw
* cell instance $456 r0 *1 8.225,17.94
X$456 89 90 91 27 92 30 257 258 cell_2rw
* cell instance $457 r0 *1 9.4,17.94
X$457 93 94 95 27 96 30 257 258 cell_2rw
* cell instance $458 r0 *1 10.575,17.94
X$458 97 98 99 27 100 30 257 258 cell_2rw
* cell instance $459 r0 *1 11.75,17.94
X$459 101 102 103 27 104 30 257 258 cell_2rw
* cell instance $460 r0 *1 12.925,17.94
X$460 105 106 107 27 108 30 257 258 cell_2rw
* cell instance $461 r0 *1 14.1,17.94
X$461 109 110 111 27 112 30 257 258 cell_2rw
* cell instance $462 r0 *1 15.275,17.94
X$462 113 114 115 27 116 30 257 258 cell_2rw
* cell instance $463 r0 *1 16.45,17.94
X$463 117 118 119 27 120 30 257 258 cell_2rw
* cell instance $464 r0 *1 17.625,17.94
X$464 121 122 123 27 124 30 257 258 cell_2rw
* cell instance $465 r0 *1 18.8,17.94
X$465 129 130 131 27 132 30 257 258 cell_2rw
* cell instance $466 r0 *1 19.975,17.94
X$466 133 134 135 27 136 30 257 258 cell_2rw
* cell instance $467 r0 *1 21.15,17.94
X$467 137 138 139 27 140 30 257 258 cell_2rw
* cell instance $468 r0 *1 22.325,17.94
X$468 141 142 143 27 144 30 257 258 cell_2rw
* cell instance $469 r0 *1 23.5,17.94
X$469 145 146 147 27 148 30 257 258 cell_2rw
* cell instance $470 r0 *1 24.675,17.94
X$470 149 150 151 27 152 30 257 258 cell_2rw
* cell instance $471 r0 *1 25.85,17.94
X$471 153 154 155 27 156 30 257 258 cell_2rw
* cell instance $472 r0 *1 27.025,17.94
X$472 157 158 159 27 160 30 257 258 cell_2rw
* cell instance $473 r0 *1 28.2,17.94
X$473 161 162 163 27 164 30 257 258 cell_2rw
* cell instance $474 r0 *1 29.375,17.94
X$474 165 166 167 27 168 30 257 258 cell_2rw
* cell instance $475 r0 *1 30.55,17.94
X$475 169 170 171 27 172 30 257 258 cell_2rw
* cell instance $476 r0 *1 31.725,17.94
X$476 173 174 175 27 176 30 257 258 cell_2rw
* cell instance $477 r0 *1 32.9,17.94
X$477 177 178 179 27 180 30 257 258 cell_2rw
* cell instance $478 r0 *1 34.075,17.94
X$478 181 182 183 27 184 30 257 258 cell_2rw
* cell instance $479 r0 *1 35.25,17.94
X$479 185 186 187 27 188 30 257 258 cell_2rw
* cell instance $480 r0 *1 36.425,17.94
X$480 189 190 191 27 192 30 257 258 cell_2rw
* cell instance $481 r0 *1 1.175,23.92
X$481 65 66 67 31 68 33 257 258 cell_2rw
* cell instance $482 r0 *1 0,23.92
X$482 61 62 63 31 64 33 257 258 cell_2rw
* cell instance $483 r0 *1 2.35,23.92
X$483 69 70 71 31 72 33 257 258 cell_2rw
* cell instance $484 r0 *1 3.525,23.92
X$484 73 74 75 31 76 33 257 258 cell_2rw
* cell instance $485 r0 *1 4.7,23.92
X$485 77 78 79 31 80 33 257 258 cell_2rw
* cell instance $486 r0 *1 5.875,23.92
X$486 81 82 83 31 84 33 257 258 cell_2rw
* cell instance $487 r0 *1 7.05,23.92
X$487 85 86 87 31 88 33 257 258 cell_2rw
* cell instance $488 r0 *1 8.225,23.92
X$488 89 90 91 31 92 33 257 258 cell_2rw
* cell instance $489 r0 *1 9.4,23.92
X$489 93 94 95 31 96 33 257 258 cell_2rw
* cell instance $490 r0 *1 10.575,23.92
X$490 97 98 99 31 100 33 257 258 cell_2rw
* cell instance $491 r0 *1 11.75,23.92
X$491 101 102 103 31 104 33 257 258 cell_2rw
* cell instance $492 r0 *1 12.925,23.92
X$492 105 106 107 31 108 33 257 258 cell_2rw
* cell instance $493 r0 *1 14.1,23.92
X$493 109 110 111 31 112 33 257 258 cell_2rw
* cell instance $494 r0 *1 15.275,23.92
X$494 113 114 115 31 116 33 257 258 cell_2rw
* cell instance $495 r0 *1 16.45,23.92
X$495 117 118 119 31 120 33 257 258 cell_2rw
* cell instance $496 r0 *1 17.625,23.92
X$496 121 122 123 31 124 33 257 258 cell_2rw
* cell instance $497 r0 *1 18.8,23.92
X$497 129 130 131 31 132 33 257 258 cell_2rw
* cell instance $498 r0 *1 19.975,23.92
X$498 133 134 135 31 136 33 257 258 cell_2rw
* cell instance $499 r0 *1 21.15,23.92
X$499 137 138 139 31 140 33 257 258 cell_2rw
* cell instance $500 r0 *1 22.325,23.92
X$500 141 142 143 31 144 33 257 258 cell_2rw
* cell instance $501 r0 *1 23.5,23.92
X$501 145 146 147 31 148 33 257 258 cell_2rw
* cell instance $502 r0 *1 24.675,23.92
X$502 149 150 151 31 152 33 257 258 cell_2rw
* cell instance $503 r0 *1 25.85,23.92
X$503 153 154 155 31 156 33 257 258 cell_2rw
* cell instance $504 r0 *1 27.025,23.92
X$504 157 158 159 31 160 33 257 258 cell_2rw
* cell instance $505 r0 *1 28.2,23.92
X$505 161 162 163 31 164 33 257 258 cell_2rw
* cell instance $506 r0 *1 29.375,23.92
X$506 165 166 167 31 168 33 257 258 cell_2rw
* cell instance $507 r0 *1 30.55,23.92
X$507 169 170 171 31 172 33 257 258 cell_2rw
* cell instance $508 r0 *1 31.725,23.92
X$508 173 174 175 31 176 33 257 258 cell_2rw
* cell instance $509 r0 *1 32.9,23.92
X$509 177 178 179 31 180 33 257 258 cell_2rw
* cell instance $510 r0 *1 34.075,23.92
X$510 181 182 183 31 184 33 257 258 cell_2rw
* cell instance $511 r0 *1 35.25,23.92
X$511 185 186 187 31 188 33 257 258 cell_2rw
* cell instance $512 r0 *1 36.425,23.92
X$512 189 190 191 31 192 33 257 258 cell_2rw
* cell instance $513 m0 *1 1.175,26.91
X$513 65 66 67 34 68 32 257 258 cell_2rw
* cell instance $514 m0 *1 0,26.91
X$514 61 62 63 34 64 32 257 258 cell_2rw
* cell instance $515 m0 *1 2.35,26.91
X$515 69 70 71 34 72 32 257 258 cell_2rw
* cell instance $516 m0 *1 3.525,26.91
X$516 73 74 75 34 76 32 257 258 cell_2rw
* cell instance $517 m0 *1 4.7,26.91
X$517 77 78 79 34 80 32 257 258 cell_2rw
* cell instance $518 m0 *1 5.875,26.91
X$518 81 82 83 34 84 32 257 258 cell_2rw
* cell instance $519 m0 *1 7.05,26.91
X$519 85 86 87 34 88 32 257 258 cell_2rw
* cell instance $520 m0 *1 8.225,26.91
X$520 89 90 91 34 92 32 257 258 cell_2rw
* cell instance $521 m0 *1 9.4,26.91
X$521 93 94 95 34 96 32 257 258 cell_2rw
* cell instance $522 m0 *1 10.575,26.91
X$522 97 98 99 34 100 32 257 258 cell_2rw
* cell instance $523 m0 *1 11.75,26.91
X$523 101 102 103 34 104 32 257 258 cell_2rw
* cell instance $524 m0 *1 12.925,26.91
X$524 105 106 107 34 108 32 257 258 cell_2rw
* cell instance $525 m0 *1 14.1,26.91
X$525 109 110 111 34 112 32 257 258 cell_2rw
* cell instance $526 m0 *1 15.275,26.91
X$526 113 114 115 34 116 32 257 258 cell_2rw
* cell instance $527 m0 *1 16.45,26.91
X$527 117 118 119 34 120 32 257 258 cell_2rw
* cell instance $528 m0 *1 17.625,26.91
X$528 121 122 123 34 124 32 257 258 cell_2rw
* cell instance $529 m0 *1 18.8,26.91
X$529 129 130 131 34 132 32 257 258 cell_2rw
* cell instance $530 m0 *1 19.975,26.91
X$530 133 134 135 34 136 32 257 258 cell_2rw
* cell instance $531 m0 *1 21.15,26.91
X$531 137 138 139 34 140 32 257 258 cell_2rw
* cell instance $532 m0 *1 22.325,26.91
X$532 141 142 143 34 144 32 257 258 cell_2rw
* cell instance $533 m0 *1 23.5,26.91
X$533 145 146 147 34 148 32 257 258 cell_2rw
* cell instance $534 m0 *1 24.675,26.91
X$534 149 150 151 34 152 32 257 258 cell_2rw
* cell instance $535 m0 *1 25.85,26.91
X$535 153 154 155 34 156 32 257 258 cell_2rw
* cell instance $536 m0 *1 27.025,26.91
X$536 157 158 159 34 160 32 257 258 cell_2rw
* cell instance $537 m0 *1 28.2,26.91
X$537 161 162 163 34 164 32 257 258 cell_2rw
* cell instance $538 m0 *1 29.375,26.91
X$538 165 166 167 34 168 32 257 258 cell_2rw
* cell instance $539 m0 *1 30.55,26.91
X$539 169 170 171 34 172 32 257 258 cell_2rw
* cell instance $540 m0 *1 31.725,26.91
X$540 173 174 175 34 176 32 257 258 cell_2rw
* cell instance $541 m0 *1 32.9,26.91
X$541 177 178 179 34 180 32 257 258 cell_2rw
* cell instance $542 m0 *1 34.075,26.91
X$542 181 182 183 34 184 32 257 258 cell_2rw
* cell instance $543 m0 *1 35.25,26.91
X$543 185 186 187 34 188 32 257 258 cell_2rw
* cell instance $544 m0 *1 36.425,26.91
X$544 189 190 191 34 192 32 257 258 cell_2rw
* cell instance $545 m0 *1 1.175,23.92
X$545 65 66 67 35 68 36 257 258 cell_2rw
* cell instance $546 m0 *1 0,23.92
X$546 61 62 63 35 64 36 257 258 cell_2rw
* cell instance $547 m0 *1 2.35,23.92
X$547 69 70 71 35 72 36 257 258 cell_2rw
* cell instance $548 m0 *1 3.525,23.92
X$548 73 74 75 35 76 36 257 258 cell_2rw
* cell instance $549 m0 *1 4.7,23.92
X$549 77 78 79 35 80 36 257 258 cell_2rw
* cell instance $550 m0 *1 5.875,23.92
X$550 81 82 83 35 84 36 257 258 cell_2rw
* cell instance $551 m0 *1 7.05,23.92
X$551 85 86 87 35 88 36 257 258 cell_2rw
* cell instance $552 m0 *1 8.225,23.92
X$552 89 90 91 35 92 36 257 258 cell_2rw
* cell instance $553 m0 *1 9.4,23.92
X$553 93 94 95 35 96 36 257 258 cell_2rw
* cell instance $554 m0 *1 10.575,23.92
X$554 97 98 99 35 100 36 257 258 cell_2rw
* cell instance $555 m0 *1 11.75,23.92
X$555 101 102 103 35 104 36 257 258 cell_2rw
* cell instance $556 m0 *1 12.925,23.92
X$556 105 106 107 35 108 36 257 258 cell_2rw
* cell instance $557 m0 *1 14.1,23.92
X$557 109 110 111 35 112 36 257 258 cell_2rw
* cell instance $558 m0 *1 15.275,23.92
X$558 113 114 115 35 116 36 257 258 cell_2rw
* cell instance $559 m0 *1 16.45,23.92
X$559 117 118 119 35 120 36 257 258 cell_2rw
* cell instance $560 m0 *1 17.625,23.92
X$560 121 122 123 35 124 36 257 258 cell_2rw
* cell instance $561 m0 *1 18.8,23.92
X$561 129 130 131 35 132 36 257 258 cell_2rw
* cell instance $562 m0 *1 19.975,23.92
X$562 133 134 135 35 136 36 257 258 cell_2rw
* cell instance $563 m0 *1 21.15,23.92
X$563 137 138 139 35 140 36 257 258 cell_2rw
* cell instance $564 m0 *1 22.325,23.92
X$564 141 142 143 35 144 36 257 258 cell_2rw
* cell instance $565 m0 *1 23.5,23.92
X$565 145 146 147 35 148 36 257 258 cell_2rw
* cell instance $566 m0 *1 24.675,23.92
X$566 149 150 151 35 152 36 257 258 cell_2rw
* cell instance $567 m0 *1 25.85,23.92
X$567 153 154 155 35 156 36 257 258 cell_2rw
* cell instance $568 m0 *1 27.025,23.92
X$568 157 158 159 35 160 36 257 258 cell_2rw
* cell instance $569 m0 *1 28.2,23.92
X$569 161 162 163 35 164 36 257 258 cell_2rw
* cell instance $570 m0 *1 29.375,23.92
X$570 165 166 167 35 168 36 257 258 cell_2rw
* cell instance $571 m0 *1 30.55,23.92
X$571 169 170 171 35 172 36 257 258 cell_2rw
* cell instance $572 m0 *1 31.725,23.92
X$572 173 174 175 35 176 36 257 258 cell_2rw
* cell instance $573 m0 *1 32.9,23.92
X$573 177 178 179 35 180 36 257 258 cell_2rw
* cell instance $574 m0 *1 34.075,23.92
X$574 181 182 183 35 184 36 257 258 cell_2rw
* cell instance $575 m0 *1 35.25,23.92
X$575 185 186 187 35 188 36 257 258 cell_2rw
* cell instance $576 m0 *1 36.425,23.92
X$576 189 190 191 35 192 36 257 258 cell_2rw
* cell instance $577 r0 *1 1.175,29.9
X$577 65 66 67 37 68 38 257 258 cell_2rw
* cell instance $578 r0 *1 0,29.9
X$578 61 62 63 37 64 38 257 258 cell_2rw
* cell instance $579 r0 *1 2.35,29.9
X$579 69 70 71 37 72 38 257 258 cell_2rw
* cell instance $580 r0 *1 3.525,29.9
X$580 73 74 75 37 76 38 257 258 cell_2rw
* cell instance $581 r0 *1 4.7,29.9
X$581 77 78 79 37 80 38 257 258 cell_2rw
* cell instance $582 r0 *1 5.875,29.9
X$582 81 82 83 37 84 38 257 258 cell_2rw
* cell instance $583 r0 *1 7.05,29.9
X$583 85 86 87 37 88 38 257 258 cell_2rw
* cell instance $584 r0 *1 8.225,29.9
X$584 89 90 91 37 92 38 257 258 cell_2rw
* cell instance $585 r0 *1 9.4,29.9
X$585 93 94 95 37 96 38 257 258 cell_2rw
* cell instance $586 r0 *1 10.575,29.9
X$586 97 98 99 37 100 38 257 258 cell_2rw
* cell instance $587 r0 *1 11.75,29.9
X$587 101 102 103 37 104 38 257 258 cell_2rw
* cell instance $588 r0 *1 12.925,29.9
X$588 105 106 107 37 108 38 257 258 cell_2rw
* cell instance $589 r0 *1 14.1,29.9
X$589 109 110 111 37 112 38 257 258 cell_2rw
* cell instance $590 r0 *1 15.275,29.9
X$590 113 114 115 37 116 38 257 258 cell_2rw
* cell instance $591 r0 *1 16.45,29.9
X$591 117 118 119 37 120 38 257 258 cell_2rw
* cell instance $592 r0 *1 17.625,29.9
X$592 121 122 123 37 124 38 257 258 cell_2rw
* cell instance $593 r0 *1 18.8,29.9
X$593 129 130 131 37 132 38 257 258 cell_2rw
* cell instance $594 r0 *1 19.975,29.9
X$594 133 134 135 37 136 38 257 258 cell_2rw
* cell instance $595 r0 *1 21.15,29.9
X$595 137 138 139 37 140 38 257 258 cell_2rw
* cell instance $596 r0 *1 22.325,29.9
X$596 141 142 143 37 144 38 257 258 cell_2rw
* cell instance $597 r0 *1 23.5,29.9
X$597 145 146 147 37 148 38 257 258 cell_2rw
* cell instance $598 r0 *1 24.675,29.9
X$598 149 150 151 37 152 38 257 258 cell_2rw
* cell instance $599 r0 *1 25.85,29.9
X$599 153 154 155 37 156 38 257 258 cell_2rw
* cell instance $600 r0 *1 27.025,29.9
X$600 157 158 159 37 160 38 257 258 cell_2rw
* cell instance $601 r0 *1 28.2,29.9
X$601 161 162 163 37 164 38 257 258 cell_2rw
* cell instance $602 r0 *1 29.375,29.9
X$602 165 166 167 37 168 38 257 258 cell_2rw
* cell instance $603 r0 *1 30.55,29.9
X$603 169 170 171 37 172 38 257 258 cell_2rw
* cell instance $604 r0 *1 31.725,29.9
X$604 173 174 175 37 176 38 257 258 cell_2rw
* cell instance $605 r0 *1 32.9,29.9
X$605 177 178 179 37 180 38 257 258 cell_2rw
* cell instance $606 r0 *1 34.075,29.9
X$606 181 182 183 37 184 38 257 258 cell_2rw
* cell instance $607 r0 *1 35.25,29.9
X$607 185 186 187 37 188 38 257 258 cell_2rw
* cell instance $608 r0 *1 36.425,29.9
X$608 189 190 191 37 192 38 257 258 cell_2rw
* cell instance $609 r0 *1 1.175,26.91
X$609 65 66 67 42 68 39 257 258 cell_2rw
* cell instance $610 r0 *1 0,26.91
X$610 61 62 63 42 64 39 257 258 cell_2rw
* cell instance $611 r0 *1 2.35,26.91
X$611 69 70 71 42 72 39 257 258 cell_2rw
* cell instance $612 r0 *1 3.525,26.91
X$612 73 74 75 42 76 39 257 258 cell_2rw
* cell instance $613 r0 *1 4.7,26.91
X$613 77 78 79 42 80 39 257 258 cell_2rw
* cell instance $614 r0 *1 5.875,26.91
X$614 81 82 83 42 84 39 257 258 cell_2rw
* cell instance $615 r0 *1 7.05,26.91
X$615 85 86 87 42 88 39 257 258 cell_2rw
* cell instance $616 r0 *1 8.225,26.91
X$616 89 90 91 42 92 39 257 258 cell_2rw
* cell instance $617 r0 *1 9.4,26.91
X$617 93 94 95 42 96 39 257 258 cell_2rw
* cell instance $618 r0 *1 10.575,26.91
X$618 97 98 99 42 100 39 257 258 cell_2rw
* cell instance $619 r0 *1 11.75,26.91
X$619 101 102 103 42 104 39 257 258 cell_2rw
* cell instance $620 r0 *1 12.925,26.91
X$620 105 106 107 42 108 39 257 258 cell_2rw
* cell instance $621 r0 *1 14.1,26.91
X$621 109 110 111 42 112 39 257 258 cell_2rw
* cell instance $622 r0 *1 15.275,26.91
X$622 113 114 115 42 116 39 257 258 cell_2rw
* cell instance $623 r0 *1 16.45,26.91
X$623 117 118 119 42 120 39 257 258 cell_2rw
* cell instance $624 r0 *1 17.625,26.91
X$624 121 122 123 42 124 39 257 258 cell_2rw
* cell instance $625 r0 *1 18.8,26.91
X$625 129 130 131 42 132 39 257 258 cell_2rw
* cell instance $626 r0 *1 19.975,26.91
X$626 133 134 135 42 136 39 257 258 cell_2rw
* cell instance $627 r0 *1 21.15,26.91
X$627 137 138 139 42 140 39 257 258 cell_2rw
* cell instance $628 r0 *1 22.325,26.91
X$628 141 142 143 42 144 39 257 258 cell_2rw
* cell instance $629 r0 *1 23.5,26.91
X$629 145 146 147 42 148 39 257 258 cell_2rw
* cell instance $630 r0 *1 24.675,26.91
X$630 149 150 151 42 152 39 257 258 cell_2rw
* cell instance $631 r0 *1 25.85,26.91
X$631 153 154 155 42 156 39 257 258 cell_2rw
* cell instance $632 r0 *1 27.025,26.91
X$632 157 158 159 42 160 39 257 258 cell_2rw
* cell instance $633 r0 *1 28.2,26.91
X$633 161 162 163 42 164 39 257 258 cell_2rw
* cell instance $634 r0 *1 29.375,26.91
X$634 165 166 167 42 168 39 257 258 cell_2rw
* cell instance $635 r0 *1 30.55,26.91
X$635 169 170 171 42 172 39 257 258 cell_2rw
* cell instance $636 r0 *1 31.725,26.91
X$636 173 174 175 42 176 39 257 258 cell_2rw
* cell instance $637 r0 *1 32.9,26.91
X$637 177 178 179 42 180 39 257 258 cell_2rw
* cell instance $638 r0 *1 34.075,26.91
X$638 181 182 183 42 184 39 257 258 cell_2rw
* cell instance $639 r0 *1 35.25,26.91
X$639 185 186 187 42 188 39 257 258 cell_2rw
* cell instance $640 r0 *1 36.425,26.91
X$640 189 190 191 42 192 39 257 258 cell_2rw
* cell instance $641 m0 *1 1.175,29.9
X$641 65 66 67 41 68 40 257 258 cell_2rw
* cell instance $642 m0 *1 0,29.9
X$642 61 62 63 41 64 40 257 258 cell_2rw
* cell instance $643 m0 *1 2.35,29.9
X$643 69 70 71 41 72 40 257 258 cell_2rw
* cell instance $644 m0 *1 3.525,29.9
X$644 73 74 75 41 76 40 257 258 cell_2rw
* cell instance $645 m0 *1 4.7,29.9
X$645 77 78 79 41 80 40 257 258 cell_2rw
* cell instance $646 m0 *1 5.875,29.9
X$646 81 82 83 41 84 40 257 258 cell_2rw
* cell instance $647 m0 *1 7.05,29.9
X$647 85 86 87 41 88 40 257 258 cell_2rw
* cell instance $648 m0 *1 8.225,29.9
X$648 89 90 91 41 92 40 257 258 cell_2rw
* cell instance $649 m0 *1 9.4,29.9
X$649 93 94 95 41 96 40 257 258 cell_2rw
* cell instance $650 m0 *1 10.575,29.9
X$650 97 98 99 41 100 40 257 258 cell_2rw
* cell instance $651 m0 *1 11.75,29.9
X$651 101 102 103 41 104 40 257 258 cell_2rw
* cell instance $652 m0 *1 12.925,29.9
X$652 105 106 107 41 108 40 257 258 cell_2rw
* cell instance $653 m0 *1 14.1,29.9
X$653 109 110 111 41 112 40 257 258 cell_2rw
* cell instance $654 m0 *1 15.275,29.9
X$654 113 114 115 41 116 40 257 258 cell_2rw
* cell instance $655 m0 *1 16.45,29.9
X$655 117 118 119 41 120 40 257 258 cell_2rw
* cell instance $656 m0 *1 17.625,29.9
X$656 121 122 123 41 124 40 257 258 cell_2rw
* cell instance $657 m0 *1 18.8,29.9
X$657 129 130 131 41 132 40 257 258 cell_2rw
* cell instance $658 m0 *1 19.975,29.9
X$658 133 134 135 41 136 40 257 258 cell_2rw
* cell instance $659 m0 *1 21.15,29.9
X$659 137 138 139 41 140 40 257 258 cell_2rw
* cell instance $660 m0 *1 22.325,29.9
X$660 141 142 143 41 144 40 257 258 cell_2rw
* cell instance $661 m0 *1 23.5,29.9
X$661 145 146 147 41 148 40 257 258 cell_2rw
* cell instance $662 m0 *1 24.675,29.9
X$662 149 150 151 41 152 40 257 258 cell_2rw
* cell instance $663 m0 *1 25.85,29.9
X$663 153 154 155 41 156 40 257 258 cell_2rw
* cell instance $664 m0 *1 27.025,29.9
X$664 157 158 159 41 160 40 257 258 cell_2rw
* cell instance $665 m0 *1 28.2,29.9
X$665 161 162 163 41 164 40 257 258 cell_2rw
* cell instance $666 m0 *1 29.375,29.9
X$666 165 166 167 41 168 40 257 258 cell_2rw
* cell instance $667 m0 *1 30.55,29.9
X$667 169 170 171 41 172 40 257 258 cell_2rw
* cell instance $668 m0 *1 31.725,29.9
X$668 173 174 175 41 176 40 257 258 cell_2rw
* cell instance $669 m0 *1 32.9,29.9
X$669 177 178 179 41 180 40 257 258 cell_2rw
* cell instance $670 m0 *1 34.075,29.9
X$670 181 182 183 41 184 40 257 258 cell_2rw
* cell instance $671 m0 *1 35.25,29.9
X$671 185 186 187 41 188 40 257 258 cell_2rw
* cell instance $672 m0 *1 36.425,29.9
X$672 189 190 191 41 192 40 257 258 cell_2rw
* cell instance $673 r0 *1 1.175,32.89
X$673 65 66 67 44 68 43 257 258 cell_2rw
* cell instance $674 r0 *1 0,32.89
X$674 61 62 63 44 64 43 257 258 cell_2rw
* cell instance $675 r0 *1 2.35,32.89
X$675 69 70 71 44 72 43 257 258 cell_2rw
* cell instance $676 r0 *1 3.525,32.89
X$676 73 74 75 44 76 43 257 258 cell_2rw
* cell instance $677 r0 *1 4.7,32.89
X$677 77 78 79 44 80 43 257 258 cell_2rw
* cell instance $678 r0 *1 5.875,32.89
X$678 81 82 83 44 84 43 257 258 cell_2rw
* cell instance $679 r0 *1 7.05,32.89
X$679 85 86 87 44 88 43 257 258 cell_2rw
* cell instance $680 r0 *1 8.225,32.89
X$680 89 90 91 44 92 43 257 258 cell_2rw
* cell instance $681 r0 *1 9.4,32.89
X$681 93 94 95 44 96 43 257 258 cell_2rw
* cell instance $682 r0 *1 10.575,32.89
X$682 97 98 99 44 100 43 257 258 cell_2rw
* cell instance $683 r0 *1 11.75,32.89
X$683 101 102 103 44 104 43 257 258 cell_2rw
* cell instance $684 r0 *1 12.925,32.89
X$684 105 106 107 44 108 43 257 258 cell_2rw
* cell instance $685 r0 *1 14.1,32.89
X$685 109 110 111 44 112 43 257 258 cell_2rw
* cell instance $686 r0 *1 15.275,32.89
X$686 113 114 115 44 116 43 257 258 cell_2rw
* cell instance $687 r0 *1 16.45,32.89
X$687 117 118 119 44 120 43 257 258 cell_2rw
* cell instance $688 r0 *1 17.625,32.89
X$688 121 122 123 44 124 43 257 258 cell_2rw
* cell instance $689 r0 *1 18.8,32.89
X$689 129 130 131 44 132 43 257 258 cell_2rw
* cell instance $690 r0 *1 19.975,32.89
X$690 133 134 135 44 136 43 257 258 cell_2rw
* cell instance $691 r0 *1 21.15,32.89
X$691 137 138 139 44 140 43 257 258 cell_2rw
* cell instance $692 r0 *1 22.325,32.89
X$692 141 142 143 44 144 43 257 258 cell_2rw
* cell instance $693 r0 *1 23.5,32.89
X$693 145 146 147 44 148 43 257 258 cell_2rw
* cell instance $694 r0 *1 24.675,32.89
X$694 149 150 151 44 152 43 257 258 cell_2rw
* cell instance $695 r0 *1 25.85,32.89
X$695 153 154 155 44 156 43 257 258 cell_2rw
* cell instance $696 r0 *1 27.025,32.89
X$696 157 158 159 44 160 43 257 258 cell_2rw
* cell instance $697 r0 *1 28.2,32.89
X$697 161 162 163 44 164 43 257 258 cell_2rw
* cell instance $698 r0 *1 29.375,32.89
X$698 165 166 167 44 168 43 257 258 cell_2rw
* cell instance $699 r0 *1 30.55,32.89
X$699 169 170 171 44 172 43 257 258 cell_2rw
* cell instance $700 r0 *1 31.725,32.89
X$700 173 174 175 44 176 43 257 258 cell_2rw
* cell instance $701 r0 *1 32.9,32.89
X$701 177 178 179 44 180 43 257 258 cell_2rw
* cell instance $702 r0 *1 34.075,32.89
X$702 181 182 183 44 184 43 257 258 cell_2rw
* cell instance $703 r0 *1 35.25,32.89
X$703 185 186 187 44 188 43 257 258 cell_2rw
* cell instance $704 r0 *1 36.425,32.89
X$704 189 190 191 44 192 43 257 258 cell_2rw
* cell instance $705 m0 *1 1.175,35.88
X$705 65 66 67 45 68 46 257 258 cell_2rw
* cell instance $706 m0 *1 0,35.88
X$706 61 62 63 45 64 46 257 258 cell_2rw
* cell instance $707 m0 *1 2.35,35.88
X$707 69 70 71 45 72 46 257 258 cell_2rw
* cell instance $708 m0 *1 3.525,35.88
X$708 73 74 75 45 76 46 257 258 cell_2rw
* cell instance $709 m0 *1 4.7,35.88
X$709 77 78 79 45 80 46 257 258 cell_2rw
* cell instance $710 m0 *1 5.875,35.88
X$710 81 82 83 45 84 46 257 258 cell_2rw
* cell instance $711 m0 *1 7.05,35.88
X$711 85 86 87 45 88 46 257 258 cell_2rw
* cell instance $712 m0 *1 8.225,35.88
X$712 89 90 91 45 92 46 257 258 cell_2rw
* cell instance $713 m0 *1 9.4,35.88
X$713 93 94 95 45 96 46 257 258 cell_2rw
* cell instance $714 m0 *1 10.575,35.88
X$714 97 98 99 45 100 46 257 258 cell_2rw
* cell instance $715 m0 *1 11.75,35.88
X$715 101 102 103 45 104 46 257 258 cell_2rw
* cell instance $716 m0 *1 12.925,35.88
X$716 105 106 107 45 108 46 257 258 cell_2rw
* cell instance $717 m0 *1 14.1,35.88
X$717 109 110 111 45 112 46 257 258 cell_2rw
* cell instance $718 m0 *1 15.275,35.88
X$718 113 114 115 45 116 46 257 258 cell_2rw
* cell instance $719 m0 *1 16.45,35.88
X$719 117 118 119 45 120 46 257 258 cell_2rw
* cell instance $720 m0 *1 17.625,35.88
X$720 121 122 123 45 124 46 257 258 cell_2rw
* cell instance $721 m0 *1 18.8,35.88
X$721 129 130 131 45 132 46 257 258 cell_2rw
* cell instance $722 m0 *1 19.975,35.88
X$722 133 134 135 45 136 46 257 258 cell_2rw
* cell instance $723 m0 *1 21.15,35.88
X$723 137 138 139 45 140 46 257 258 cell_2rw
* cell instance $724 m0 *1 22.325,35.88
X$724 141 142 143 45 144 46 257 258 cell_2rw
* cell instance $725 m0 *1 23.5,35.88
X$725 145 146 147 45 148 46 257 258 cell_2rw
* cell instance $726 m0 *1 24.675,35.88
X$726 149 150 151 45 152 46 257 258 cell_2rw
* cell instance $727 m0 *1 25.85,35.88
X$727 153 154 155 45 156 46 257 258 cell_2rw
* cell instance $728 m0 *1 27.025,35.88
X$728 157 158 159 45 160 46 257 258 cell_2rw
* cell instance $729 m0 *1 28.2,35.88
X$729 161 162 163 45 164 46 257 258 cell_2rw
* cell instance $730 m0 *1 29.375,35.88
X$730 165 166 167 45 168 46 257 258 cell_2rw
* cell instance $731 m0 *1 30.55,35.88
X$731 169 170 171 45 172 46 257 258 cell_2rw
* cell instance $732 m0 *1 31.725,35.88
X$732 173 174 175 45 176 46 257 258 cell_2rw
* cell instance $733 m0 *1 32.9,35.88
X$733 177 178 179 45 180 46 257 258 cell_2rw
* cell instance $734 m0 *1 34.075,35.88
X$734 181 182 183 45 184 46 257 258 cell_2rw
* cell instance $735 m0 *1 35.25,35.88
X$735 185 186 187 45 188 46 257 258 cell_2rw
* cell instance $736 m0 *1 36.425,35.88
X$736 189 190 191 45 192 46 257 258 cell_2rw
* cell instance $737 m0 *1 1.175,32.89
X$737 65 66 67 48 68 47 257 258 cell_2rw
* cell instance $738 m0 *1 0,32.89
X$738 61 62 63 48 64 47 257 258 cell_2rw
* cell instance $739 m0 *1 2.35,32.89
X$739 69 70 71 48 72 47 257 258 cell_2rw
* cell instance $740 m0 *1 3.525,32.89
X$740 73 74 75 48 76 47 257 258 cell_2rw
* cell instance $741 m0 *1 4.7,32.89
X$741 77 78 79 48 80 47 257 258 cell_2rw
* cell instance $742 m0 *1 5.875,32.89
X$742 81 82 83 48 84 47 257 258 cell_2rw
* cell instance $743 m0 *1 7.05,32.89
X$743 85 86 87 48 88 47 257 258 cell_2rw
* cell instance $744 m0 *1 8.225,32.89
X$744 89 90 91 48 92 47 257 258 cell_2rw
* cell instance $745 m0 *1 9.4,32.89
X$745 93 94 95 48 96 47 257 258 cell_2rw
* cell instance $746 m0 *1 10.575,32.89
X$746 97 98 99 48 100 47 257 258 cell_2rw
* cell instance $747 m0 *1 11.75,32.89
X$747 101 102 103 48 104 47 257 258 cell_2rw
* cell instance $748 m0 *1 12.925,32.89
X$748 105 106 107 48 108 47 257 258 cell_2rw
* cell instance $749 m0 *1 14.1,32.89
X$749 109 110 111 48 112 47 257 258 cell_2rw
* cell instance $750 m0 *1 15.275,32.89
X$750 113 114 115 48 116 47 257 258 cell_2rw
* cell instance $751 m0 *1 16.45,32.89
X$751 117 118 119 48 120 47 257 258 cell_2rw
* cell instance $752 m0 *1 17.625,32.89
X$752 121 122 123 48 124 47 257 258 cell_2rw
* cell instance $753 m0 *1 18.8,32.89
X$753 129 130 131 48 132 47 257 258 cell_2rw
* cell instance $754 m0 *1 19.975,32.89
X$754 133 134 135 48 136 47 257 258 cell_2rw
* cell instance $755 m0 *1 21.15,32.89
X$755 137 138 139 48 140 47 257 258 cell_2rw
* cell instance $756 m0 *1 22.325,32.89
X$756 141 142 143 48 144 47 257 258 cell_2rw
* cell instance $757 m0 *1 23.5,32.89
X$757 145 146 147 48 148 47 257 258 cell_2rw
* cell instance $758 m0 *1 24.675,32.89
X$758 149 150 151 48 152 47 257 258 cell_2rw
* cell instance $759 m0 *1 25.85,32.89
X$759 153 154 155 48 156 47 257 258 cell_2rw
* cell instance $760 m0 *1 27.025,32.89
X$760 157 158 159 48 160 47 257 258 cell_2rw
* cell instance $761 m0 *1 28.2,32.89
X$761 161 162 163 48 164 47 257 258 cell_2rw
* cell instance $762 m0 *1 29.375,32.89
X$762 165 166 167 48 168 47 257 258 cell_2rw
* cell instance $763 m0 *1 30.55,32.89
X$763 169 170 171 48 172 47 257 258 cell_2rw
* cell instance $764 m0 *1 31.725,32.89
X$764 173 174 175 48 176 47 257 258 cell_2rw
* cell instance $765 m0 *1 32.9,32.89
X$765 177 178 179 48 180 47 257 258 cell_2rw
* cell instance $766 m0 *1 34.075,32.89
X$766 181 182 183 48 184 47 257 258 cell_2rw
* cell instance $767 m0 *1 35.25,32.89
X$767 185 186 187 48 188 47 257 258 cell_2rw
* cell instance $768 m0 *1 36.425,32.89
X$768 189 190 191 48 192 47 257 258 cell_2rw
* cell instance $769 m0 *1 1.175,38.87
X$769 65 66 67 54 68 49 257 258 cell_2rw
* cell instance $770 m0 *1 0,38.87
X$770 61 62 63 54 64 49 257 258 cell_2rw
* cell instance $771 m0 *1 2.35,38.87
X$771 69 70 71 54 72 49 257 258 cell_2rw
* cell instance $772 m0 *1 3.525,38.87
X$772 73 74 75 54 76 49 257 258 cell_2rw
* cell instance $773 m0 *1 4.7,38.87
X$773 77 78 79 54 80 49 257 258 cell_2rw
* cell instance $774 m0 *1 5.875,38.87
X$774 81 82 83 54 84 49 257 258 cell_2rw
* cell instance $775 m0 *1 7.05,38.87
X$775 85 86 87 54 88 49 257 258 cell_2rw
* cell instance $776 m0 *1 8.225,38.87
X$776 89 90 91 54 92 49 257 258 cell_2rw
* cell instance $777 m0 *1 9.4,38.87
X$777 93 94 95 54 96 49 257 258 cell_2rw
* cell instance $778 m0 *1 10.575,38.87
X$778 97 98 99 54 100 49 257 258 cell_2rw
* cell instance $779 m0 *1 11.75,38.87
X$779 101 102 103 54 104 49 257 258 cell_2rw
* cell instance $780 m0 *1 12.925,38.87
X$780 105 106 107 54 108 49 257 258 cell_2rw
* cell instance $781 m0 *1 14.1,38.87
X$781 109 110 111 54 112 49 257 258 cell_2rw
* cell instance $782 m0 *1 15.275,38.87
X$782 113 114 115 54 116 49 257 258 cell_2rw
* cell instance $783 m0 *1 16.45,38.87
X$783 117 118 119 54 120 49 257 258 cell_2rw
* cell instance $784 m0 *1 17.625,38.87
X$784 121 122 123 54 124 49 257 258 cell_2rw
* cell instance $785 m0 *1 18.8,38.87
X$785 129 130 131 54 132 49 257 258 cell_2rw
* cell instance $786 m0 *1 19.975,38.87
X$786 133 134 135 54 136 49 257 258 cell_2rw
* cell instance $787 m0 *1 21.15,38.87
X$787 137 138 139 54 140 49 257 258 cell_2rw
* cell instance $788 m0 *1 22.325,38.87
X$788 141 142 143 54 144 49 257 258 cell_2rw
* cell instance $789 m0 *1 23.5,38.87
X$789 145 146 147 54 148 49 257 258 cell_2rw
* cell instance $790 m0 *1 24.675,38.87
X$790 149 150 151 54 152 49 257 258 cell_2rw
* cell instance $791 m0 *1 25.85,38.87
X$791 153 154 155 54 156 49 257 258 cell_2rw
* cell instance $792 m0 *1 27.025,38.87
X$792 157 158 159 54 160 49 257 258 cell_2rw
* cell instance $793 m0 *1 28.2,38.87
X$793 161 162 163 54 164 49 257 258 cell_2rw
* cell instance $794 m0 *1 29.375,38.87
X$794 165 166 167 54 168 49 257 258 cell_2rw
* cell instance $795 m0 *1 30.55,38.87
X$795 169 170 171 54 172 49 257 258 cell_2rw
* cell instance $796 m0 *1 31.725,38.87
X$796 173 174 175 54 176 49 257 258 cell_2rw
* cell instance $797 m0 *1 32.9,38.87
X$797 177 178 179 54 180 49 257 258 cell_2rw
* cell instance $798 m0 *1 34.075,38.87
X$798 181 182 183 54 184 49 257 258 cell_2rw
* cell instance $799 m0 *1 35.25,38.87
X$799 185 186 187 54 188 49 257 258 cell_2rw
* cell instance $800 m0 *1 36.425,38.87
X$800 189 190 191 54 192 49 257 258 cell_2rw
* cell instance $801 r0 *1 1.175,38.87
X$801 65 66 67 51 68 50 257 258 cell_2rw
* cell instance $802 r0 *1 0,38.87
X$802 61 62 63 51 64 50 257 258 cell_2rw
* cell instance $803 r0 *1 2.35,38.87
X$803 69 70 71 51 72 50 257 258 cell_2rw
* cell instance $804 r0 *1 3.525,38.87
X$804 73 74 75 51 76 50 257 258 cell_2rw
* cell instance $805 r0 *1 4.7,38.87
X$805 77 78 79 51 80 50 257 258 cell_2rw
* cell instance $806 r0 *1 5.875,38.87
X$806 81 82 83 51 84 50 257 258 cell_2rw
* cell instance $807 r0 *1 7.05,38.87
X$807 85 86 87 51 88 50 257 258 cell_2rw
* cell instance $808 r0 *1 8.225,38.87
X$808 89 90 91 51 92 50 257 258 cell_2rw
* cell instance $809 r0 *1 9.4,38.87
X$809 93 94 95 51 96 50 257 258 cell_2rw
* cell instance $810 r0 *1 10.575,38.87
X$810 97 98 99 51 100 50 257 258 cell_2rw
* cell instance $811 r0 *1 11.75,38.87
X$811 101 102 103 51 104 50 257 258 cell_2rw
* cell instance $812 r0 *1 12.925,38.87
X$812 105 106 107 51 108 50 257 258 cell_2rw
* cell instance $813 r0 *1 14.1,38.87
X$813 109 110 111 51 112 50 257 258 cell_2rw
* cell instance $814 r0 *1 15.275,38.87
X$814 113 114 115 51 116 50 257 258 cell_2rw
* cell instance $815 r0 *1 16.45,38.87
X$815 117 118 119 51 120 50 257 258 cell_2rw
* cell instance $816 r0 *1 17.625,38.87
X$816 121 122 123 51 124 50 257 258 cell_2rw
* cell instance $817 r0 *1 18.8,38.87
X$817 129 130 131 51 132 50 257 258 cell_2rw
* cell instance $818 r0 *1 19.975,38.87
X$818 133 134 135 51 136 50 257 258 cell_2rw
* cell instance $819 r0 *1 21.15,38.87
X$819 137 138 139 51 140 50 257 258 cell_2rw
* cell instance $820 r0 *1 22.325,38.87
X$820 141 142 143 51 144 50 257 258 cell_2rw
* cell instance $821 r0 *1 23.5,38.87
X$821 145 146 147 51 148 50 257 258 cell_2rw
* cell instance $822 r0 *1 24.675,38.87
X$822 149 150 151 51 152 50 257 258 cell_2rw
* cell instance $823 r0 *1 25.85,38.87
X$823 153 154 155 51 156 50 257 258 cell_2rw
* cell instance $824 r0 *1 27.025,38.87
X$824 157 158 159 51 160 50 257 258 cell_2rw
* cell instance $825 r0 *1 28.2,38.87
X$825 161 162 163 51 164 50 257 258 cell_2rw
* cell instance $826 r0 *1 29.375,38.87
X$826 165 166 167 51 168 50 257 258 cell_2rw
* cell instance $827 r0 *1 30.55,38.87
X$827 169 170 171 51 172 50 257 258 cell_2rw
* cell instance $828 r0 *1 31.725,38.87
X$828 173 174 175 51 176 50 257 258 cell_2rw
* cell instance $829 r0 *1 32.9,38.87
X$829 177 178 179 51 180 50 257 258 cell_2rw
* cell instance $830 r0 *1 34.075,38.87
X$830 181 182 183 51 184 50 257 258 cell_2rw
* cell instance $831 r0 *1 35.25,38.87
X$831 185 186 187 51 188 50 257 258 cell_2rw
* cell instance $832 r0 *1 36.425,38.87
X$832 189 190 191 51 192 50 257 258 cell_2rw
* cell instance $833 r0 *1 1.175,35.88
X$833 65 66 67 53 68 52 257 258 cell_2rw
* cell instance $834 r0 *1 0,35.88
X$834 61 62 63 53 64 52 257 258 cell_2rw
* cell instance $835 r0 *1 2.35,35.88
X$835 69 70 71 53 72 52 257 258 cell_2rw
* cell instance $836 r0 *1 3.525,35.88
X$836 73 74 75 53 76 52 257 258 cell_2rw
* cell instance $837 r0 *1 4.7,35.88
X$837 77 78 79 53 80 52 257 258 cell_2rw
* cell instance $838 r0 *1 5.875,35.88
X$838 81 82 83 53 84 52 257 258 cell_2rw
* cell instance $839 r0 *1 7.05,35.88
X$839 85 86 87 53 88 52 257 258 cell_2rw
* cell instance $840 r0 *1 8.225,35.88
X$840 89 90 91 53 92 52 257 258 cell_2rw
* cell instance $841 r0 *1 9.4,35.88
X$841 93 94 95 53 96 52 257 258 cell_2rw
* cell instance $842 r0 *1 10.575,35.88
X$842 97 98 99 53 100 52 257 258 cell_2rw
* cell instance $843 r0 *1 11.75,35.88
X$843 101 102 103 53 104 52 257 258 cell_2rw
* cell instance $844 r0 *1 12.925,35.88
X$844 105 106 107 53 108 52 257 258 cell_2rw
* cell instance $845 r0 *1 14.1,35.88
X$845 109 110 111 53 112 52 257 258 cell_2rw
* cell instance $846 r0 *1 15.275,35.88
X$846 113 114 115 53 116 52 257 258 cell_2rw
* cell instance $847 r0 *1 16.45,35.88
X$847 117 118 119 53 120 52 257 258 cell_2rw
* cell instance $848 r0 *1 17.625,35.88
X$848 121 122 123 53 124 52 257 258 cell_2rw
* cell instance $849 r0 *1 18.8,35.88
X$849 129 130 131 53 132 52 257 258 cell_2rw
* cell instance $850 r0 *1 19.975,35.88
X$850 133 134 135 53 136 52 257 258 cell_2rw
* cell instance $851 r0 *1 21.15,35.88
X$851 137 138 139 53 140 52 257 258 cell_2rw
* cell instance $852 r0 *1 22.325,35.88
X$852 141 142 143 53 144 52 257 258 cell_2rw
* cell instance $853 r0 *1 23.5,35.88
X$853 145 146 147 53 148 52 257 258 cell_2rw
* cell instance $854 r0 *1 24.675,35.88
X$854 149 150 151 53 152 52 257 258 cell_2rw
* cell instance $855 r0 *1 25.85,35.88
X$855 153 154 155 53 156 52 257 258 cell_2rw
* cell instance $856 r0 *1 27.025,35.88
X$856 157 158 159 53 160 52 257 258 cell_2rw
* cell instance $857 r0 *1 28.2,35.88
X$857 161 162 163 53 164 52 257 258 cell_2rw
* cell instance $858 r0 *1 29.375,35.88
X$858 165 166 167 53 168 52 257 258 cell_2rw
* cell instance $859 r0 *1 30.55,35.88
X$859 169 170 171 53 172 52 257 258 cell_2rw
* cell instance $860 r0 *1 31.725,35.88
X$860 173 174 175 53 176 52 257 258 cell_2rw
* cell instance $861 r0 *1 32.9,35.88
X$861 177 178 179 53 180 52 257 258 cell_2rw
* cell instance $862 r0 *1 34.075,35.88
X$862 181 182 183 53 184 52 257 258 cell_2rw
* cell instance $863 r0 *1 35.25,35.88
X$863 185 186 187 53 188 52 257 258 cell_2rw
* cell instance $864 r0 *1 36.425,35.88
X$864 189 190 191 53 192 52 257 258 cell_2rw
* cell instance $865 r0 *1 1.175,41.86
X$865 65 66 67 56 68 55 257 258 cell_2rw
* cell instance $866 r0 *1 0,41.86
X$866 61 62 63 56 64 55 257 258 cell_2rw
* cell instance $867 r0 *1 2.35,41.86
X$867 69 70 71 56 72 55 257 258 cell_2rw
* cell instance $868 r0 *1 3.525,41.86
X$868 73 74 75 56 76 55 257 258 cell_2rw
* cell instance $869 r0 *1 4.7,41.86
X$869 77 78 79 56 80 55 257 258 cell_2rw
* cell instance $870 r0 *1 5.875,41.86
X$870 81 82 83 56 84 55 257 258 cell_2rw
* cell instance $871 r0 *1 7.05,41.86
X$871 85 86 87 56 88 55 257 258 cell_2rw
* cell instance $872 r0 *1 8.225,41.86
X$872 89 90 91 56 92 55 257 258 cell_2rw
* cell instance $873 r0 *1 9.4,41.86
X$873 93 94 95 56 96 55 257 258 cell_2rw
* cell instance $874 r0 *1 10.575,41.86
X$874 97 98 99 56 100 55 257 258 cell_2rw
* cell instance $875 r0 *1 11.75,41.86
X$875 101 102 103 56 104 55 257 258 cell_2rw
* cell instance $876 r0 *1 12.925,41.86
X$876 105 106 107 56 108 55 257 258 cell_2rw
* cell instance $877 r0 *1 14.1,41.86
X$877 109 110 111 56 112 55 257 258 cell_2rw
* cell instance $878 r0 *1 15.275,41.86
X$878 113 114 115 56 116 55 257 258 cell_2rw
* cell instance $879 r0 *1 16.45,41.86
X$879 117 118 119 56 120 55 257 258 cell_2rw
* cell instance $880 r0 *1 17.625,41.86
X$880 121 122 123 56 124 55 257 258 cell_2rw
* cell instance $881 r0 *1 18.8,41.86
X$881 129 130 131 56 132 55 257 258 cell_2rw
* cell instance $882 r0 *1 19.975,41.86
X$882 133 134 135 56 136 55 257 258 cell_2rw
* cell instance $883 r0 *1 21.15,41.86
X$883 137 138 139 56 140 55 257 258 cell_2rw
* cell instance $884 r0 *1 22.325,41.86
X$884 141 142 143 56 144 55 257 258 cell_2rw
* cell instance $885 r0 *1 23.5,41.86
X$885 145 146 147 56 148 55 257 258 cell_2rw
* cell instance $886 r0 *1 24.675,41.86
X$886 149 150 151 56 152 55 257 258 cell_2rw
* cell instance $887 r0 *1 25.85,41.86
X$887 153 154 155 56 156 55 257 258 cell_2rw
* cell instance $888 r0 *1 27.025,41.86
X$888 157 158 159 56 160 55 257 258 cell_2rw
* cell instance $889 r0 *1 28.2,41.86
X$889 161 162 163 56 164 55 257 258 cell_2rw
* cell instance $890 r0 *1 29.375,41.86
X$890 165 166 167 56 168 55 257 258 cell_2rw
* cell instance $891 r0 *1 30.55,41.86
X$891 169 170 171 56 172 55 257 258 cell_2rw
* cell instance $892 r0 *1 31.725,41.86
X$892 173 174 175 56 176 55 257 258 cell_2rw
* cell instance $893 r0 *1 32.9,41.86
X$893 177 178 179 56 180 55 257 258 cell_2rw
* cell instance $894 r0 *1 34.075,41.86
X$894 181 182 183 56 184 55 257 258 cell_2rw
* cell instance $895 r0 *1 35.25,41.86
X$895 185 186 187 56 188 55 257 258 cell_2rw
* cell instance $896 r0 *1 36.425,41.86
X$896 189 190 191 56 192 55 257 258 cell_2rw
* cell instance $897 m0 *1 1.175,44.85
X$897 65 66 67 60 68 57 257 258 cell_2rw
* cell instance $898 m0 *1 0,44.85
X$898 61 62 63 60 64 57 257 258 cell_2rw
* cell instance $899 m0 *1 2.35,44.85
X$899 69 70 71 60 72 57 257 258 cell_2rw
* cell instance $900 m0 *1 3.525,44.85
X$900 73 74 75 60 76 57 257 258 cell_2rw
* cell instance $901 m0 *1 4.7,44.85
X$901 77 78 79 60 80 57 257 258 cell_2rw
* cell instance $902 m0 *1 5.875,44.85
X$902 81 82 83 60 84 57 257 258 cell_2rw
* cell instance $903 m0 *1 7.05,44.85
X$903 85 86 87 60 88 57 257 258 cell_2rw
* cell instance $904 m0 *1 8.225,44.85
X$904 89 90 91 60 92 57 257 258 cell_2rw
* cell instance $905 m0 *1 9.4,44.85
X$905 93 94 95 60 96 57 257 258 cell_2rw
* cell instance $906 m0 *1 10.575,44.85
X$906 97 98 99 60 100 57 257 258 cell_2rw
* cell instance $907 m0 *1 11.75,44.85
X$907 101 102 103 60 104 57 257 258 cell_2rw
* cell instance $908 m0 *1 12.925,44.85
X$908 105 106 107 60 108 57 257 258 cell_2rw
* cell instance $909 m0 *1 14.1,44.85
X$909 109 110 111 60 112 57 257 258 cell_2rw
* cell instance $910 m0 *1 15.275,44.85
X$910 113 114 115 60 116 57 257 258 cell_2rw
* cell instance $911 m0 *1 16.45,44.85
X$911 117 118 119 60 120 57 257 258 cell_2rw
* cell instance $912 m0 *1 17.625,44.85
X$912 121 122 123 60 124 57 257 258 cell_2rw
* cell instance $913 m0 *1 18.8,44.85
X$913 129 130 131 60 132 57 257 258 cell_2rw
* cell instance $914 m0 *1 19.975,44.85
X$914 133 134 135 60 136 57 257 258 cell_2rw
* cell instance $915 m0 *1 21.15,44.85
X$915 137 138 139 60 140 57 257 258 cell_2rw
* cell instance $916 m0 *1 22.325,44.85
X$916 141 142 143 60 144 57 257 258 cell_2rw
* cell instance $917 m0 *1 23.5,44.85
X$917 145 146 147 60 148 57 257 258 cell_2rw
* cell instance $918 m0 *1 24.675,44.85
X$918 149 150 151 60 152 57 257 258 cell_2rw
* cell instance $919 m0 *1 25.85,44.85
X$919 153 154 155 60 156 57 257 258 cell_2rw
* cell instance $920 m0 *1 27.025,44.85
X$920 157 158 159 60 160 57 257 258 cell_2rw
* cell instance $921 m0 *1 28.2,44.85
X$921 161 162 163 60 164 57 257 258 cell_2rw
* cell instance $922 m0 *1 29.375,44.85
X$922 165 166 167 60 168 57 257 258 cell_2rw
* cell instance $923 m0 *1 30.55,44.85
X$923 169 170 171 60 172 57 257 258 cell_2rw
* cell instance $924 m0 *1 31.725,44.85
X$924 173 174 175 60 176 57 257 258 cell_2rw
* cell instance $925 m0 *1 32.9,44.85
X$925 177 178 179 60 180 57 257 258 cell_2rw
* cell instance $926 m0 *1 34.075,44.85
X$926 181 182 183 60 184 57 257 258 cell_2rw
* cell instance $927 m0 *1 35.25,44.85
X$927 185 186 187 60 188 57 257 258 cell_2rw
* cell instance $928 m0 *1 36.425,44.85
X$928 189 190 191 60 192 57 257 258 cell_2rw
* cell instance $929 m0 *1 1.175,41.86
X$929 65 66 67 59 68 58 257 258 cell_2rw
* cell instance $930 m0 *1 0,41.86
X$930 61 62 63 59 64 58 257 258 cell_2rw
* cell instance $931 m0 *1 2.35,41.86
X$931 69 70 71 59 72 58 257 258 cell_2rw
* cell instance $932 m0 *1 3.525,41.86
X$932 73 74 75 59 76 58 257 258 cell_2rw
* cell instance $933 m0 *1 4.7,41.86
X$933 77 78 79 59 80 58 257 258 cell_2rw
* cell instance $934 m0 *1 5.875,41.86
X$934 81 82 83 59 84 58 257 258 cell_2rw
* cell instance $935 m0 *1 7.05,41.86
X$935 85 86 87 59 88 58 257 258 cell_2rw
* cell instance $936 m0 *1 8.225,41.86
X$936 89 90 91 59 92 58 257 258 cell_2rw
* cell instance $937 m0 *1 9.4,41.86
X$937 93 94 95 59 96 58 257 258 cell_2rw
* cell instance $938 m0 *1 10.575,41.86
X$938 97 98 99 59 100 58 257 258 cell_2rw
* cell instance $939 m0 *1 11.75,41.86
X$939 101 102 103 59 104 58 257 258 cell_2rw
* cell instance $940 m0 *1 12.925,41.86
X$940 105 106 107 59 108 58 257 258 cell_2rw
* cell instance $941 m0 *1 14.1,41.86
X$941 109 110 111 59 112 58 257 258 cell_2rw
* cell instance $942 m0 *1 15.275,41.86
X$942 113 114 115 59 116 58 257 258 cell_2rw
* cell instance $943 m0 *1 16.45,41.86
X$943 117 118 119 59 120 58 257 258 cell_2rw
* cell instance $944 m0 *1 17.625,41.86
X$944 121 122 123 59 124 58 257 258 cell_2rw
* cell instance $945 m0 *1 18.8,41.86
X$945 129 130 131 59 132 58 257 258 cell_2rw
* cell instance $946 m0 *1 19.975,41.86
X$946 133 134 135 59 136 58 257 258 cell_2rw
* cell instance $947 m0 *1 21.15,41.86
X$947 137 138 139 59 140 58 257 258 cell_2rw
* cell instance $948 m0 *1 22.325,41.86
X$948 141 142 143 59 144 58 257 258 cell_2rw
* cell instance $949 m0 *1 23.5,41.86
X$949 145 146 147 59 148 58 257 258 cell_2rw
* cell instance $950 m0 *1 24.675,41.86
X$950 149 150 151 59 152 58 257 258 cell_2rw
* cell instance $951 m0 *1 25.85,41.86
X$951 153 154 155 59 156 58 257 258 cell_2rw
* cell instance $952 m0 *1 27.025,41.86
X$952 157 158 159 59 160 58 257 258 cell_2rw
* cell instance $953 m0 *1 28.2,41.86
X$953 161 162 163 59 164 58 257 258 cell_2rw
* cell instance $954 m0 *1 29.375,41.86
X$954 165 166 167 59 168 58 257 258 cell_2rw
* cell instance $955 m0 *1 30.55,41.86
X$955 169 170 171 59 172 58 257 258 cell_2rw
* cell instance $956 m0 *1 31.725,41.86
X$956 173 174 175 59 176 58 257 258 cell_2rw
* cell instance $957 m0 *1 32.9,41.86
X$957 177 178 179 59 180 58 257 258 cell_2rw
* cell instance $958 m0 *1 34.075,41.86
X$958 181 182 183 59 184 58 257 258 cell_2rw
* cell instance $959 m0 *1 35.25,41.86
X$959 185 186 187 59 188 58 257 258 cell_2rw
* cell instance $960 m0 *1 36.425,41.86
X$960 189 190 191 59 192 58 257 258 cell_2rw
* cell instance $961 r0 *1 0,44.85
X$961 61 62 63 127 64 128 257 258 cell_2rw
* cell instance $962 m0 *1 0,47.84
X$962 61 62 63 126 64 125 257 258 cell_2rw
* cell instance $963 m0 *1 0,50.83
X$963 61 62 63 195 64 197 257 258 cell_2rw
* cell instance $964 r0 *1 0,47.84
X$964 61 62 63 199 64 201 257 258 cell_2rw
* cell instance $965 r0 *1 0,50.83
X$965 61 62 63 202 64 194 257 258 cell_2rw
* cell instance $966 m0 *1 0,53.82
X$966 61 62 63 198 64 193 257 258 cell_2rw
* cell instance $967 r0 *1 0,53.82
X$967 61 62 63 196 64 200 257 258 cell_2rw
* cell instance $968 m0 *1 0,56.81
X$968 61 62 63 203 64 207 257 258 cell_2rw
* cell instance $969 r0 *1 0,56.81
X$969 61 62 63 206 64 208 257 258 cell_2rw
* cell instance $970 m0 *1 0,59.8
X$970 61 62 63 205 64 204 257 258 cell_2rw
* cell instance $971 r0 *1 0,59.8
X$971 61 62 63 214 64 213 257 258 cell_2rw
* cell instance $972 m0 *1 0,62.79
X$972 61 62 63 212 64 211 257 258 cell_2rw
* cell instance $973 r0 *1 0,62.79
X$973 61 62 63 210 64 209 257 258 cell_2rw
* cell instance $974 m0 *1 0,65.78
X$974 61 62 63 219 64 217 257 258 cell_2rw
* cell instance $975 r0 *1 0,65.78
X$975 61 62 63 216 64 215 257 258 cell_2rw
* cell instance $976 m0 *1 0,68.77
X$976 61 62 63 218 64 220 257 258 cell_2rw
* cell instance $977 r0 *1 0,68.77
X$977 61 62 63 224 64 223 257 258 cell_2rw
* cell instance $978 m0 *1 0,71.76
X$978 61 62 63 221 64 222 257 258 cell_2rw
* cell instance $979 r0 *1 0,71.76
X$979 61 62 63 226 64 225 257 258 cell_2rw
* cell instance $980 m0 *1 0,74.75
X$980 61 62 63 231 64 232 257 258 cell_2rw
* cell instance $981 r0 *1 0,74.75
X$981 61 62 63 230 64 229 257 258 cell_2rw
* cell instance $982 m0 *1 0,77.74
X$982 61 62 63 227 64 228 257 258 cell_2rw
* cell instance $983 m0 *1 0,80.73
X$983 61 62 63 233 64 236 257 258 cell_2rw
* cell instance $984 r0 *1 0,77.74
X$984 61 62 63 237 64 238 257 258 cell_2rw
* cell instance $985 r0 *1 0,80.73
X$985 61 62 63 235 64 234 257 258 cell_2rw
* cell instance $986 m0 *1 0,83.72
X$986 61 62 63 240 64 242 257 258 cell_2rw
* cell instance $987 m0 *1 0,86.71
X$987 61 62 63 244 64 243 257 258 cell_2rw
* cell instance $988 r0 *1 0,83.72
X$988 61 62 63 239 64 241 257 258 cell_2rw
* cell instance $989 r0 *1 0,86.71
X$989 61 62 63 245 64 247 257 258 cell_2rw
* cell instance $990 m0 *1 0,89.7
X$990 61 62 63 250 64 249 257 258 cell_2rw
* cell instance $991 r0 *1 0,89.7
X$991 61 62 63 246 64 248 257 258 cell_2rw
* cell instance $992 m0 *1 0,92.69
X$992 61 62 63 253 64 256 257 258 cell_2rw
* cell instance $993 r0 *1 0,92.69
X$993 61 62 63 255 64 254 257 258 cell_2rw
* cell instance $994 m0 *1 0,95.68
X$994 61 62 63 251 64 252 257 258 cell_2rw
* cell instance $995 r0 *1 1.175,44.85
X$995 65 66 67 127 68 128 257 258 cell_2rw
* cell instance $996 m0 *1 1.175,47.84
X$996 65 66 67 126 68 125 257 258 cell_2rw
* cell instance $997 m0 *1 1.175,50.83
X$997 65 66 67 195 68 197 257 258 cell_2rw
* cell instance $998 r0 *1 1.175,47.84
X$998 65 66 67 199 68 201 257 258 cell_2rw
* cell instance $999 r0 *1 1.175,50.83
X$999 65 66 67 202 68 194 257 258 cell_2rw
* cell instance $1000 m0 *1 1.175,53.82
X$1000 65 66 67 198 68 193 257 258 cell_2rw
* cell instance $1001 r0 *1 1.175,53.82
X$1001 65 66 67 196 68 200 257 258 cell_2rw
* cell instance $1002 m0 *1 1.175,56.81
X$1002 65 66 67 203 68 207 257 258 cell_2rw
* cell instance $1003 r0 *1 1.175,56.81
X$1003 65 66 67 206 68 208 257 258 cell_2rw
* cell instance $1004 m0 *1 1.175,59.8
X$1004 65 66 67 205 68 204 257 258 cell_2rw
* cell instance $1005 r0 *1 1.175,59.8
X$1005 65 66 67 214 68 213 257 258 cell_2rw
* cell instance $1006 m0 *1 1.175,62.79
X$1006 65 66 67 212 68 211 257 258 cell_2rw
* cell instance $1007 r0 *1 1.175,62.79
X$1007 65 66 67 210 68 209 257 258 cell_2rw
* cell instance $1008 m0 *1 1.175,65.78
X$1008 65 66 67 219 68 217 257 258 cell_2rw
* cell instance $1009 r0 *1 1.175,65.78
X$1009 65 66 67 216 68 215 257 258 cell_2rw
* cell instance $1010 m0 *1 1.175,68.77
X$1010 65 66 67 218 68 220 257 258 cell_2rw
* cell instance $1011 r0 *1 1.175,68.77
X$1011 65 66 67 224 68 223 257 258 cell_2rw
* cell instance $1012 m0 *1 1.175,71.76
X$1012 65 66 67 221 68 222 257 258 cell_2rw
* cell instance $1013 r0 *1 1.175,71.76
X$1013 65 66 67 226 68 225 257 258 cell_2rw
* cell instance $1014 m0 *1 1.175,74.75
X$1014 65 66 67 231 68 232 257 258 cell_2rw
* cell instance $1015 r0 *1 1.175,74.75
X$1015 65 66 67 230 68 229 257 258 cell_2rw
* cell instance $1016 m0 *1 1.175,77.74
X$1016 65 66 67 227 68 228 257 258 cell_2rw
* cell instance $1017 r0 *1 1.175,77.74
X$1017 65 66 67 237 68 238 257 258 cell_2rw
* cell instance $1018 m0 *1 1.175,80.73
X$1018 65 66 67 233 68 236 257 258 cell_2rw
* cell instance $1019 m0 *1 1.175,83.72
X$1019 65 66 67 240 68 242 257 258 cell_2rw
* cell instance $1020 r0 *1 1.175,80.73
X$1020 65 66 67 235 68 234 257 258 cell_2rw
* cell instance $1021 r0 *1 1.175,83.72
X$1021 65 66 67 239 68 241 257 258 cell_2rw
* cell instance $1022 m0 *1 1.175,86.71
X$1022 65 66 67 244 68 243 257 258 cell_2rw
* cell instance $1023 r0 *1 1.175,86.71
X$1023 65 66 67 245 68 247 257 258 cell_2rw
* cell instance $1024 m0 *1 1.175,89.7
X$1024 65 66 67 250 68 249 257 258 cell_2rw
* cell instance $1025 r0 *1 1.175,89.7
X$1025 65 66 67 246 68 248 257 258 cell_2rw
* cell instance $1026 m0 *1 1.175,92.69
X$1026 65 66 67 253 68 256 257 258 cell_2rw
* cell instance $1027 r0 *1 1.175,92.69
X$1027 65 66 67 255 68 254 257 258 cell_2rw
* cell instance $1028 m0 *1 1.175,95.68
X$1028 65 66 67 251 68 252 257 258 cell_2rw
* cell instance $1029 m0 *1 2.35,47.84
X$1029 69 70 71 126 72 125 257 258 cell_2rw
* cell instance $1030 r0 *1 2.35,44.85
X$1030 69 70 71 127 72 128 257 258 cell_2rw
* cell instance $1031 r0 *1 2.35,47.84
X$1031 69 70 71 199 72 201 257 258 cell_2rw
* cell instance $1032 m0 *1 2.35,50.83
X$1032 69 70 71 195 72 197 257 258 cell_2rw
* cell instance $1033 r0 *1 2.35,50.83
X$1033 69 70 71 202 72 194 257 258 cell_2rw
* cell instance $1034 m0 *1 2.35,53.82
X$1034 69 70 71 198 72 193 257 258 cell_2rw
* cell instance $1035 m0 *1 2.35,56.81
X$1035 69 70 71 203 72 207 257 258 cell_2rw
* cell instance $1036 r0 *1 2.35,53.82
X$1036 69 70 71 196 72 200 257 258 cell_2rw
* cell instance $1037 r0 *1 2.35,56.81
X$1037 69 70 71 206 72 208 257 258 cell_2rw
* cell instance $1038 m0 *1 2.35,59.8
X$1038 69 70 71 205 72 204 257 258 cell_2rw
* cell instance $1039 m0 *1 2.35,62.79
X$1039 69 70 71 212 72 211 257 258 cell_2rw
* cell instance $1040 r0 *1 2.35,59.8
X$1040 69 70 71 214 72 213 257 258 cell_2rw
* cell instance $1041 r0 *1 2.35,62.79
X$1041 69 70 71 210 72 209 257 258 cell_2rw
* cell instance $1042 m0 *1 2.35,65.78
X$1042 69 70 71 219 72 217 257 258 cell_2rw
* cell instance $1043 r0 *1 2.35,65.78
X$1043 69 70 71 216 72 215 257 258 cell_2rw
* cell instance $1044 m0 *1 2.35,68.77
X$1044 69 70 71 218 72 220 257 258 cell_2rw
* cell instance $1045 m0 *1 2.35,71.76
X$1045 69 70 71 221 72 222 257 258 cell_2rw
* cell instance $1046 r0 *1 2.35,68.77
X$1046 69 70 71 224 72 223 257 258 cell_2rw
* cell instance $1047 m0 *1 2.35,74.75
X$1047 69 70 71 231 72 232 257 258 cell_2rw
* cell instance $1048 r0 *1 2.35,71.76
X$1048 69 70 71 226 72 225 257 258 cell_2rw
* cell instance $1049 r0 *1 2.35,74.75
X$1049 69 70 71 230 72 229 257 258 cell_2rw
* cell instance $1050 m0 *1 2.35,77.74
X$1050 69 70 71 227 72 228 257 258 cell_2rw
* cell instance $1051 r0 *1 2.35,77.74
X$1051 69 70 71 237 72 238 257 258 cell_2rw
* cell instance $1052 m0 *1 2.35,80.73
X$1052 69 70 71 233 72 236 257 258 cell_2rw
* cell instance $1053 r0 *1 2.35,80.73
X$1053 69 70 71 235 72 234 257 258 cell_2rw
* cell instance $1054 m0 *1 2.35,83.72
X$1054 69 70 71 240 72 242 257 258 cell_2rw
* cell instance $1055 m0 *1 2.35,86.71
X$1055 69 70 71 244 72 243 257 258 cell_2rw
* cell instance $1056 r0 *1 2.35,83.72
X$1056 69 70 71 239 72 241 257 258 cell_2rw
* cell instance $1057 r0 *1 2.35,86.71
X$1057 69 70 71 245 72 247 257 258 cell_2rw
* cell instance $1058 m0 *1 2.35,89.7
X$1058 69 70 71 250 72 249 257 258 cell_2rw
* cell instance $1059 r0 *1 2.35,89.7
X$1059 69 70 71 246 72 248 257 258 cell_2rw
* cell instance $1060 m0 *1 2.35,92.69
X$1060 69 70 71 253 72 256 257 258 cell_2rw
* cell instance $1061 r0 *1 2.35,92.69
X$1061 69 70 71 255 72 254 257 258 cell_2rw
* cell instance $1062 m0 *1 2.35,95.68
X$1062 69 70 71 251 72 252 257 258 cell_2rw
* cell instance $1063 r0 *1 3.525,44.85
X$1063 73 74 75 127 76 128 257 258 cell_2rw
* cell instance $1064 m0 *1 3.525,47.84
X$1064 73 74 75 126 76 125 257 258 cell_2rw
* cell instance $1065 m0 *1 3.525,50.83
X$1065 73 74 75 195 76 197 257 258 cell_2rw
* cell instance $1066 r0 *1 3.525,47.84
X$1066 73 74 75 199 76 201 257 258 cell_2rw
* cell instance $1067 r0 *1 3.525,50.83
X$1067 73 74 75 202 76 194 257 258 cell_2rw
* cell instance $1068 m0 *1 3.525,53.82
X$1068 73 74 75 198 76 193 257 258 cell_2rw
* cell instance $1069 r0 *1 3.525,53.82
X$1069 73 74 75 196 76 200 257 258 cell_2rw
* cell instance $1070 m0 *1 3.525,56.81
X$1070 73 74 75 203 76 207 257 258 cell_2rw
* cell instance $1071 m0 *1 3.525,59.8
X$1071 73 74 75 205 76 204 257 258 cell_2rw
* cell instance $1072 r0 *1 3.525,56.81
X$1072 73 74 75 206 76 208 257 258 cell_2rw
* cell instance $1073 r0 *1 3.525,59.8
X$1073 73 74 75 214 76 213 257 258 cell_2rw
* cell instance $1074 m0 *1 3.525,62.79
X$1074 73 74 75 212 76 211 257 258 cell_2rw
* cell instance $1075 r0 *1 3.525,62.79
X$1075 73 74 75 210 76 209 257 258 cell_2rw
* cell instance $1076 m0 *1 3.525,65.78
X$1076 73 74 75 219 76 217 257 258 cell_2rw
* cell instance $1077 r0 *1 3.525,65.78
X$1077 73 74 75 216 76 215 257 258 cell_2rw
* cell instance $1078 m0 *1 3.525,68.77
X$1078 73 74 75 218 76 220 257 258 cell_2rw
* cell instance $1079 r0 *1 3.525,68.77
X$1079 73 74 75 224 76 223 257 258 cell_2rw
* cell instance $1080 m0 *1 3.525,71.76
X$1080 73 74 75 221 76 222 257 258 cell_2rw
* cell instance $1081 r0 *1 3.525,71.76
X$1081 73 74 75 226 76 225 257 258 cell_2rw
* cell instance $1082 m0 *1 3.525,74.75
X$1082 73 74 75 231 76 232 257 258 cell_2rw
* cell instance $1083 m0 *1 3.525,77.74
X$1083 73 74 75 227 76 228 257 258 cell_2rw
* cell instance $1084 r0 *1 3.525,74.75
X$1084 73 74 75 230 76 229 257 258 cell_2rw
* cell instance $1085 r0 *1 3.525,77.74
X$1085 73 74 75 237 76 238 257 258 cell_2rw
* cell instance $1086 m0 *1 3.525,80.73
X$1086 73 74 75 233 76 236 257 258 cell_2rw
* cell instance $1087 r0 *1 3.525,80.73
X$1087 73 74 75 235 76 234 257 258 cell_2rw
* cell instance $1088 m0 *1 3.525,83.72
X$1088 73 74 75 240 76 242 257 258 cell_2rw
* cell instance $1089 r0 *1 3.525,83.72
X$1089 73 74 75 239 76 241 257 258 cell_2rw
* cell instance $1090 m0 *1 3.525,86.71
X$1090 73 74 75 244 76 243 257 258 cell_2rw
* cell instance $1091 r0 *1 3.525,86.71
X$1091 73 74 75 245 76 247 257 258 cell_2rw
* cell instance $1092 m0 *1 3.525,89.7
X$1092 73 74 75 250 76 249 257 258 cell_2rw
* cell instance $1093 r0 *1 3.525,89.7
X$1093 73 74 75 246 76 248 257 258 cell_2rw
* cell instance $1094 m0 *1 3.525,92.69
X$1094 73 74 75 253 76 256 257 258 cell_2rw
* cell instance $1095 r0 *1 3.525,92.69
X$1095 73 74 75 255 76 254 257 258 cell_2rw
* cell instance $1096 m0 *1 3.525,95.68
X$1096 73 74 75 251 76 252 257 258 cell_2rw
* cell instance $1097 r0 *1 4.7,44.85
X$1097 77 78 79 127 80 128 257 258 cell_2rw
* cell instance $1098 m0 *1 4.7,47.84
X$1098 77 78 79 126 80 125 257 258 cell_2rw
* cell instance $1099 r0 *1 4.7,47.84
X$1099 77 78 79 199 80 201 257 258 cell_2rw
* cell instance $1100 m0 *1 4.7,50.83
X$1100 77 78 79 195 80 197 257 258 cell_2rw
* cell instance $1101 r0 *1 4.7,50.83
X$1101 77 78 79 202 80 194 257 258 cell_2rw
* cell instance $1102 m0 *1 4.7,53.82
X$1102 77 78 79 198 80 193 257 258 cell_2rw
* cell instance $1103 r0 *1 4.7,53.82
X$1103 77 78 79 196 80 200 257 258 cell_2rw
* cell instance $1104 m0 *1 4.7,56.81
X$1104 77 78 79 203 80 207 257 258 cell_2rw
* cell instance $1105 r0 *1 4.7,56.81
X$1105 77 78 79 206 80 208 257 258 cell_2rw
* cell instance $1106 m0 *1 4.7,59.8
X$1106 77 78 79 205 80 204 257 258 cell_2rw
* cell instance $1107 r0 *1 4.7,59.8
X$1107 77 78 79 214 80 213 257 258 cell_2rw
* cell instance $1108 m0 *1 4.7,62.79
X$1108 77 78 79 212 80 211 257 258 cell_2rw
* cell instance $1109 r0 *1 4.7,62.79
X$1109 77 78 79 210 80 209 257 258 cell_2rw
* cell instance $1110 m0 *1 4.7,65.78
X$1110 77 78 79 219 80 217 257 258 cell_2rw
* cell instance $1111 m0 *1 4.7,68.77
X$1111 77 78 79 218 80 220 257 258 cell_2rw
* cell instance $1112 r0 *1 4.7,65.78
X$1112 77 78 79 216 80 215 257 258 cell_2rw
* cell instance $1113 r0 *1 4.7,68.77
X$1113 77 78 79 224 80 223 257 258 cell_2rw
* cell instance $1114 m0 *1 4.7,71.76
X$1114 77 78 79 221 80 222 257 258 cell_2rw
* cell instance $1115 m0 *1 4.7,74.75
X$1115 77 78 79 231 80 232 257 258 cell_2rw
* cell instance $1116 r0 *1 4.7,71.76
X$1116 77 78 79 226 80 225 257 258 cell_2rw
* cell instance $1117 r0 *1 4.7,74.75
X$1117 77 78 79 230 80 229 257 258 cell_2rw
* cell instance $1118 m0 *1 4.7,77.74
X$1118 77 78 79 227 80 228 257 258 cell_2rw
* cell instance $1119 r0 *1 4.7,77.74
X$1119 77 78 79 237 80 238 257 258 cell_2rw
* cell instance $1120 m0 *1 4.7,80.73
X$1120 77 78 79 233 80 236 257 258 cell_2rw
* cell instance $1121 r0 *1 4.7,80.73
X$1121 77 78 79 235 80 234 257 258 cell_2rw
* cell instance $1122 m0 *1 4.7,83.72
X$1122 77 78 79 240 80 242 257 258 cell_2rw
* cell instance $1123 m0 *1 4.7,86.71
X$1123 77 78 79 244 80 243 257 258 cell_2rw
* cell instance $1124 r0 *1 4.7,83.72
X$1124 77 78 79 239 80 241 257 258 cell_2rw
* cell instance $1125 m0 *1 4.7,89.7
X$1125 77 78 79 250 80 249 257 258 cell_2rw
* cell instance $1126 r0 *1 4.7,86.71
X$1126 77 78 79 245 80 247 257 258 cell_2rw
* cell instance $1127 r0 *1 4.7,89.7
X$1127 77 78 79 246 80 248 257 258 cell_2rw
* cell instance $1128 m0 *1 4.7,92.69
X$1128 77 78 79 253 80 256 257 258 cell_2rw
* cell instance $1129 r0 *1 4.7,92.69
X$1129 77 78 79 255 80 254 257 258 cell_2rw
* cell instance $1130 m0 *1 4.7,95.68
X$1130 77 78 79 251 80 252 257 258 cell_2rw
* cell instance $1131 m0 *1 5.875,47.84
X$1131 81 82 83 126 84 125 257 258 cell_2rw
* cell instance $1132 r0 *1 5.875,44.85
X$1132 81 82 83 127 84 128 257 258 cell_2rw
* cell instance $1133 r0 *1 5.875,47.84
X$1133 81 82 83 199 84 201 257 258 cell_2rw
* cell instance $1134 m0 *1 5.875,50.83
X$1134 81 82 83 195 84 197 257 258 cell_2rw
* cell instance $1135 r0 *1 5.875,50.83
X$1135 81 82 83 202 84 194 257 258 cell_2rw
* cell instance $1136 m0 *1 5.875,53.82
X$1136 81 82 83 198 84 193 257 258 cell_2rw
* cell instance $1137 r0 *1 5.875,53.82
X$1137 81 82 83 196 84 200 257 258 cell_2rw
* cell instance $1138 m0 *1 5.875,56.81
X$1138 81 82 83 203 84 207 257 258 cell_2rw
* cell instance $1139 r0 *1 5.875,56.81
X$1139 81 82 83 206 84 208 257 258 cell_2rw
* cell instance $1140 m0 *1 5.875,59.8
X$1140 81 82 83 205 84 204 257 258 cell_2rw
* cell instance $1141 r0 *1 5.875,59.8
X$1141 81 82 83 214 84 213 257 258 cell_2rw
* cell instance $1142 m0 *1 5.875,62.79
X$1142 81 82 83 212 84 211 257 258 cell_2rw
* cell instance $1143 r0 *1 5.875,62.79
X$1143 81 82 83 210 84 209 257 258 cell_2rw
* cell instance $1144 m0 *1 5.875,65.78
X$1144 81 82 83 219 84 217 257 258 cell_2rw
* cell instance $1145 r0 *1 5.875,65.78
X$1145 81 82 83 216 84 215 257 258 cell_2rw
* cell instance $1146 m0 *1 5.875,68.77
X$1146 81 82 83 218 84 220 257 258 cell_2rw
* cell instance $1147 r0 *1 5.875,68.77
X$1147 81 82 83 224 84 223 257 258 cell_2rw
* cell instance $1148 m0 *1 5.875,71.76
X$1148 81 82 83 221 84 222 257 258 cell_2rw
* cell instance $1149 r0 *1 5.875,71.76
X$1149 81 82 83 226 84 225 257 258 cell_2rw
* cell instance $1150 m0 *1 5.875,74.75
X$1150 81 82 83 231 84 232 257 258 cell_2rw
* cell instance $1151 m0 *1 5.875,77.74
X$1151 81 82 83 227 84 228 257 258 cell_2rw
* cell instance $1152 r0 *1 5.875,74.75
X$1152 81 82 83 230 84 229 257 258 cell_2rw
* cell instance $1153 r0 *1 5.875,77.74
X$1153 81 82 83 237 84 238 257 258 cell_2rw
* cell instance $1154 m0 *1 5.875,80.73
X$1154 81 82 83 233 84 236 257 258 cell_2rw
* cell instance $1155 r0 *1 5.875,80.73
X$1155 81 82 83 235 84 234 257 258 cell_2rw
* cell instance $1156 m0 *1 5.875,83.72
X$1156 81 82 83 240 84 242 257 258 cell_2rw
* cell instance $1157 r0 *1 5.875,83.72
X$1157 81 82 83 239 84 241 257 258 cell_2rw
* cell instance $1158 m0 *1 5.875,86.71
X$1158 81 82 83 244 84 243 257 258 cell_2rw
* cell instance $1159 r0 *1 5.875,86.71
X$1159 81 82 83 245 84 247 257 258 cell_2rw
* cell instance $1160 m0 *1 5.875,89.7
X$1160 81 82 83 250 84 249 257 258 cell_2rw
* cell instance $1161 r0 *1 5.875,89.7
X$1161 81 82 83 246 84 248 257 258 cell_2rw
* cell instance $1162 m0 *1 5.875,92.69
X$1162 81 82 83 253 84 256 257 258 cell_2rw
* cell instance $1163 r0 *1 5.875,92.69
X$1163 81 82 83 255 84 254 257 258 cell_2rw
* cell instance $1164 m0 *1 5.875,95.68
X$1164 81 82 83 251 84 252 257 258 cell_2rw
* cell instance $1165 r0 *1 7.05,44.85
X$1165 85 86 87 127 88 128 257 258 cell_2rw
* cell instance $1166 m0 *1 7.05,47.84
X$1166 85 86 87 126 88 125 257 258 cell_2rw
* cell instance $1167 r0 *1 7.05,47.84
X$1167 85 86 87 199 88 201 257 258 cell_2rw
* cell instance $1168 m0 *1 7.05,50.83
X$1168 85 86 87 195 88 197 257 258 cell_2rw
* cell instance $1169 r0 *1 7.05,50.83
X$1169 85 86 87 202 88 194 257 258 cell_2rw
* cell instance $1170 m0 *1 7.05,53.82
X$1170 85 86 87 198 88 193 257 258 cell_2rw
* cell instance $1171 r0 *1 7.05,53.82
X$1171 85 86 87 196 88 200 257 258 cell_2rw
* cell instance $1172 m0 *1 7.05,56.81
X$1172 85 86 87 203 88 207 257 258 cell_2rw
* cell instance $1173 r0 *1 7.05,56.81
X$1173 85 86 87 206 88 208 257 258 cell_2rw
* cell instance $1174 m0 *1 7.05,59.8
X$1174 85 86 87 205 88 204 257 258 cell_2rw
* cell instance $1175 r0 *1 7.05,59.8
X$1175 85 86 87 214 88 213 257 258 cell_2rw
* cell instance $1176 m0 *1 7.05,62.79
X$1176 85 86 87 212 88 211 257 258 cell_2rw
* cell instance $1177 r0 *1 7.05,62.79
X$1177 85 86 87 210 88 209 257 258 cell_2rw
* cell instance $1178 m0 *1 7.05,65.78
X$1178 85 86 87 219 88 217 257 258 cell_2rw
* cell instance $1179 r0 *1 7.05,65.78
X$1179 85 86 87 216 88 215 257 258 cell_2rw
* cell instance $1180 m0 *1 7.05,68.77
X$1180 85 86 87 218 88 220 257 258 cell_2rw
* cell instance $1181 r0 *1 7.05,68.77
X$1181 85 86 87 224 88 223 257 258 cell_2rw
* cell instance $1182 m0 *1 7.05,71.76
X$1182 85 86 87 221 88 222 257 258 cell_2rw
* cell instance $1183 r0 *1 7.05,71.76
X$1183 85 86 87 226 88 225 257 258 cell_2rw
* cell instance $1184 m0 *1 7.05,74.75
X$1184 85 86 87 231 88 232 257 258 cell_2rw
* cell instance $1185 r0 *1 7.05,74.75
X$1185 85 86 87 230 88 229 257 258 cell_2rw
* cell instance $1186 m0 *1 7.05,77.74
X$1186 85 86 87 227 88 228 257 258 cell_2rw
* cell instance $1187 r0 *1 7.05,77.74
X$1187 85 86 87 237 88 238 257 258 cell_2rw
* cell instance $1188 m0 *1 7.05,80.73
X$1188 85 86 87 233 88 236 257 258 cell_2rw
* cell instance $1189 m0 *1 7.05,83.72
X$1189 85 86 87 240 88 242 257 258 cell_2rw
* cell instance $1190 r0 *1 7.05,80.73
X$1190 85 86 87 235 88 234 257 258 cell_2rw
* cell instance $1191 r0 *1 7.05,83.72
X$1191 85 86 87 239 88 241 257 258 cell_2rw
* cell instance $1192 m0 *1 7.05,86.71
X$1192 85 86 87 244 88 243 257 258 cell_2rw
* cell instance $1193 r0 *1 7.05,86.71
X$1193 85 86 87 245 88 247 257 258 cell_2rw
* cell instance $1194 m0 *1 7.05,89.7
X$1194 85 86 87 250 88 249 257 258 cell_2rw
* cell instance $1195 m0 *1 7.05,92.69
X$1195 85 86 87 253 88 256 257 258 cell_2rw
* cell instance $1196 r0 *1 7.05,89.7
X$1196 85 86 87 246 88 248 257 258 cell_2rw
* cell instance $1197 m0 *1 7.05,95.68
X$1197 85 86 87 251 88 252 257 258 cell_2rw
* cell instance $1198 r0 *1 7.05,92.69
X$1198 85 86 87 255 88 254 257 258 cell_2rw
* cell instance $1199 m0 *1 8.225,47.84
X$1199 89 90 91 126 92 125 257 258 cell_2rw
* cell instance $1200 r0 *1 8.225,44.85
X$1200 89 90 91 127 92 128 257 258 cell_2rw
* cell instance $1201 m0 *1 8.225,50.83
X$1201 89 90 91 195 92 197 257 258 cell_2rw
* cell instance $1202 r0 *1 8.225,47.84
X$1202 89 90 91 199 92 201 257 258 cell_2rw
* cell instance $1203 r0 *1 8.225,50.83
X$1203 89 90 91 202 92 194 257 258 cell_2rw
* cell instance $1204 m0 *1 8.225,53.82
X$1204 89 90 91 198 92 193 257 258 cell_2rw
* cell instance $1205 r0 *1 8.225,53.82
X$1205 89 90 91 196 92 200 257 258 cell_2rw
* cell instance $1206 m0 *1 8.225,56.81
X$1206 89 90 91 203 92 207 257 258 cell_2rw
* cell instance $1207 r0 *1 8.225,56.81
X$1207 89 90 91 206 92 208 257 258 cell_2rw
* cell instance $1208 m0 *1 8.225,59.8
X$1208 89 90 91 205 92 204 257 258 cell_2rw
* cell instance $1209 r0 *1 8.225,59.8
X$1209 89 90 91 214 92 213 257 258 cell_2rw
* cell instance $1210 m0 *1 8.225,62.79
X$1210 89 90 91 212 92 211 257 258 cell_2rw
* cell instance $1211 r0 *1 8.225,62.79
X$1211 89 90 91 210 92 209 257 258 cell_2rw
* cell instance $1212 m0 *1 8.225,65.78
X$1212 89 90 91 219 92 217 257 258 cell_2rw
* cell instance $1213 r0 *1 8.225,65.78
X$1213 89 90 91 216 92 215 257 258 cell_2rw
* cell instance $1214 m0 *1 8.225,68.77
X$1214 89 90 91 218 92 220 257 258 cell_2rw
* cell instance $1215 m0 *1 8.225,71.76
X$1215 89 90 91 221 92 222 257 258 cell_2rw
* cell instance $1216 r0 *1 8.225,68.77
X$1216 89 90 91 224 92 223 257 258 cell_2rw
* cell instance $1217 m0 *1 8.225,74.75
X$1217 89 90 91 231 92 232 257 258 cell_2rw
* cell instance $1218 r0 *1 8.225,71.76
X$1218 89 90 91 226 92 225 257 258 cell_2rw
* cell instance $1219 r0 *1 8.225,74.75
X$1219 89 90 91 230 92 229 257 258 cell_2rw
* cell instance $1220 m0 *1 8.225,77.74
X$1220 89 90 91 227 92 228 257 258 cell_2rw
* cell instance $1221 r0 *1 8.225,77.74
X$1221 89 90 91 237 92 238 257 258 cell_2rw
* cell instance $1222 m0 *1 8.225,80.73
X$1222 89 90 91 233 92 236 257 258 cell_2rw
* cell instance $1223 r0 *1 8.225,80.73
X$1223 89 90 91 235 92 234 257 258 cell_2rw
* cell instance $1224 m0 *1 8.225,83.72
X$1224 89 90 91 240 92 242 257 258 cell_2rw
* cell instance $1225 r0 *1 8.225,83.72
X$1225 89 90 91 239 92 241 257 258 cell_2rw
* cell instance $1226 m0 *1 8.225,86.71
X$1226 89 90 91 244 92 243 257 258 cell_2rw
* cell instance $1227 r0 *1 8.225,86.71
X$1227 89 90 91 245 92 247 257 258 cell_2rw
* cell instance $1228 m0 *1 8.225,89.7
X$1228 89 90 91 250 92 249 257 258 cell_2rw
* cell instance $1229 r0 *1 8.225,89.7
X$1229 89 90 91 246 92 248 257 258 cell_2rw
* cell instance $1230 m0 *1 8.225,92.69
X$1230 89 90 91 253 92 256 257 258 cell_2rw
* cell instance $1231 m0 *1 8.225,95.68
X$1231 89 90 91 251 92 252 257 258 cell_2rw
* cell instance $1232 r0 *1 8.225,92.69
X$1232 89 90 91 255 92 254 257 258 cell_2rw
* cell instance $1233 r0 *1 9.4,44.85
X$1233 93 94 95 127 96 128 257 258 cell_2rw
* cell instance $1234 m0 *1 9.4,47.84
X$1234 93 94 95 126 96 125 257 258 cell_2rw
* cell instance $1235 r0 *1 9.4,47.84
X$1235 93 94 95 199 96 201 257 258 cell_2rw
* cell instance $1236 m0 *1 9.4,50.83
X$1236 93 94 95 195 96 197 257 258 cell_2rw
* cell instance $1237 r0 *1 9.4,50.83
X$1237 93 94 95 202 96 194 257 258 cell_2rw
* cell instance $1238 m0 *1 9.4,53.82
X$1238 93 94 95 198 96 193 257 258 cell_2rw
* cell instance $1239 r0 *1 9.4,53.82
X$1239 93 94 95 196 96 200 257 258 cell_2rw
* cell instance $1240 m0 *1 9.4,56.81
X$1240 93 94 95 203 96 207 257 258 cell_2rw
* cell instance $1241 r0 *1 9.4,56.81
X$1241 93 94 95 206 96 208 257 258 cell_2rw
* cell instance $1242 m0 *1 9.4,59.8
X$1242 93 94 95 205 96 204 257 258 cell_2rw
* cell instance $1243 m0 *1 9.4,62.79
X$1243 93 94 95 212 96 211 257 258 cell_2rw
* cell instance $1244 r0 *1 9.4,59.8
X$1244 93 94 95 214 96 213 257 258 cell_2rw
* cell instance $1245 r0 *1 9.4,62.79
X$1245 93 94 95 210 96 209 257 258 cell_2rw
* cell instance $1246 m0 *1 9.4,65.78
X$1246 93 94 95 219 96 217 257 258 cell_2rw
* cell instance $1247 r0 *1 9.4,65.78
X$1247 93 94 95 216 96 215 257 258 cell_2rw
* cell instance $1248 m0 *1 9.4,68.77
X$1248 93 94 95 218 96 220 257 258 cell_2rw
* cell instance $1249 r0 *1 9.4,68.77
X$1249 93 94 95 224 96 223 257 258 cell_2rw
* cell instance $1250 m0 *1 9.4,71.76
X$1250 93 94 95 221 96 222 257 258 cell_2rw
* cell instance $1251 r0 *1 9.4,71.76
X$1251 93 94 95 226 96 225 257 258 cell_2rw
* cell instance $1252 m0 *1 9.4,74.75
X$1252 93 94 95 231 96 232 257 258 cell_2rw
* cell instance $1253 r0 *1 9.4,74.75
X$1253 93 94 95 230 96 229 257 258 cell_2rw
* cell instance $1254 m0 *1 9.4,77.74
X$1254 93 94 95 227 96 228 257 258 cell_2rw
* cell instance $1255 r0 *1 9.4,77.74
X$1255 93 94 95 237 96 238 257 258 cell_2rw
* cell instance $1256 m0 *1 9.4,80.73
X$1256 93 94 95 233 96 236 257 258 cell_2rw
* cell instance $1257 r0 *1 9.4,80.73
X$1257 93 94 95 235 96 234 257 258 cell_2rw
* cell instance $1258 m0 *1 9.4,83.72
X$1258 93 94 95 240 96 242 257 258 cell_2rw
* cell instance $1259 r0 *1 9.4,83.72
X$1259 93 94 95 239 96 241 257 258 cell_2rw
* cell instance $1260 m0 *1 9.4,86.71
X$1260 93 94 95 244 96 243 257 258 cell_2rw
* cell instance $1261 m0 *1 9.4,89.7
X$1261 93 94 95 250 96 249 257 258 cell_2rw
* cell instance $1262 r0 *1 9.4,86.71
X$1262 93 94 95 245 96 247 257 258 cell_2rw
* cell instance $1263 r0 *1 9.4,89.7
X$1263 93 94 95 246 96 248 257 258 cell_2rw
* cell instance $1264 m0 *1 9.4,92.69
X$1264 93 94 95 253 96 256 257 258 cell_2rw
* cell instance $1265 m0 *1 9.4,95.68
X$1265 93 94 95 251 96 252 257 258 cell_2rw
* cell instance $1266 r0 *1 9.4,92.69
X$1266 93 94 95 255 96 254 257 258 cell_2rw
* cell instance $1267 r0 *1 10.575,44.85
X$1267 97 98 99 127 100 128 257 258 cell_2rw
* cell instance $1268 m0 *1 10.575,47.84
X$1268 97 98 99 126 100 125 257 258 cell_2rw
* cell instance $1269 r0 *1 10.575,47.84
X$1269 97 98 99 199 100 201 257 258 cell_2rw
* cell instance $1270 m0 *1 10.575,50.83
X$1270 97 98 99 195 100 197 257 258 cell_2rw
* cell instance $1271 r0 *1 10.575,50.83
X$1271 97 98 99 202 100 194 257 258 cell_2rw
* cell instance $1272 m0 *1 10.575,53.82
X$1272 97 98 99 198 100 193 257 258 cell_2rw
* cell instance $1273 r0 *1 10.575,53.82
X$1273 97 98 99 196 100 200 257 258 cell_2rw
* cell instance $1274 m0 *1 10.575,56.81
X$1274 97 98 99 203 100 207 257 258 cell_2rw
* cell instance $1275 r0 *1 10.575,56.81
X$1275 97 98 99 206 100 208 257 258 cell_2rw
* cell instance $1276 m0 *1 10.575,59.8
X$1276 97 98 99 205 100 204 257 258 cell_2rw
* cell instance $1277 r0 *1 10.575,59.8
X$1277 97 98 99 214 100 213 257 258 cell_2rw
* cell instance $1278 m0 *1 10.575,62.79
X$1278 97 98 99 212 100 211 257 258 cell_2rw
* cell instance $1279 r0 *1 10.575,62.79
X$1279 97 98 99 210 100 209 257 258 cell_2rw
* cell instance $1280 m0 *1 10.575,65.78
X$1280 97 98 99 219 100 217 257 258 cell_2rw
* cell instance $1281 r0 *1 10.575,65.78
X$1281 97 98 99 216 100 215 257 258 cell_2rw
* cell instance $1282 m0 *1 10.575,68.77
X$1282 97 98 99 218 100 220 257 258 cell_2rw
* cell instance $1283 r0 *1 10.575,68.77
X$1283 97 98 99 224 100 223 257 258 cell_2rw
* cell instance $1284 m0 *1 10.575,71.76
X$1284 97 98 99 221 100 222 257 258 cell_2rw
* cell instance $1285 r0 *1 10.575,71.76
X$1285 97 98 99 226 100 225 257 258 cell_2rw
* cell instance $1286 m0 *1 10.575,74.75
X$1286 97 98 99 231 100 232 257 258 cell_2rw
* cell instance $1287 r0 *1 10.575,74.75
X$1287 97 98 99 230 100 229 257 258 cell_2rw
* cell instance $1288 m0 *1 10.575,77.74
X$1288 97 98 99 227 100 228 257 258 cell_2rw
* cell instance $1289 r0 *1 10.575,77.74
X$1289 97 98 99 237 100 238 257 258 cell_2rw
* cell instance $1290 m0 *1 10.575,80.73
X$1290 97 98 99 233 100 236 257 258 cell_2rw
* cell instance $1291 r0 *1 10.575,80.73
X$1291 97 98 99 235 100 234 257 258 cell_2rw
* cell instance $1292 m0 *1 10.575,83.72
X$1292 97 98 99 240 100 242 257 258 cell_2rw
* cell instance $1293 m0 *1 10.575,86.71
X$1293 97 98 99 244 100 243 257 258 cell_2rw
* cell instance $1294 r0 *1 10.575,83.72
X$1294 97 98 99 239 100 241 257 258 cell_2rw
* cell instance $1295 r0 *1 10.575,86.71
X$1295 97 98 99 245 100 247 257 258 cell_2rw
* cell instance $1296 m0 *1 10.575,89.7
X$1296 97 98 99 250 100 249 257 258 cell_2rw
* cell instance $1297 r0 *1 10.575,89.7
X$1297 97 98 99 246 100 248 257 258 cell_2rw
* cell instance $1298 m0 *1 10.575,92.69
X$1298 97 98 99 253 100 256 257 258 cell_2rw
* cell instance $1299 m0 *1 10.575,95.68
X$1299 97 98 99 251 100 252 257 258 cell_2rw
* cell instance $1300 r0 *1 10.575,92.69
X$1300 97 98 99 255 100 254 257 258 cell_2rw
* cell instance $1301 m0 *1 11.75,47.84
X$1301 101 102 103 126 104 125 257 258 cell_2rw
* cell instance $1302 r0 *1 11.75,44.85
X$1302 101 102 103 127 104 128 257 258 cell_2rw
* cell instance $1303 r0 *1 11.75,47.84
X$1303 101 102 103 199 104 201 257 258 cell_2rw
* cell instance $1304 m0 *1 11.75,50.83
X$1304 101 102 103 195 104 197 257 258 cell_2rw
* cell instance $1305 m0 *1 11.75,53.82
X$1305 101 102 103 198 104 193 257 258 cell_2rw
* cell instance $1306 r0 *1 11.75,50.83
X$1306 101 102 103 202 104 194 257 258 cell_2rw
* cell instance $1307 r0 *1 11.75,53.82
X$1307 101 102 103 196 104 200 257 258 cell_2rw
* cell instance $1308 m0 *1 11.75,56.81
X$1308 101 102 103 203 104 207 257 258 cell_2rw
* cell instance $1309 r0 *1 11.75,56.81
X$1309 101 102 103 206 104 208 257 258 cell_2rw
* cell instance $1310 m0 *1 11.75,59.8
X$1310 101 102 103 205 104 204 257 258 cell_2rw
* cell instance $1311 r0 *1 11.75,59.8
X$1311 101 102 103 214 104 213 257 258 cell_2rw
* cell instance $1312 m0 *1 11.75,62.79
X$1312 101 102 103 212 104 211 257 258 cell_2rw
* cell instance $1313 m0 *1 11.75,65.78
X$1313 101 102 103 219 104 217 257 258 cell_2rw
* cell instance $1314 r0 *1 11.75,62.79
X$1314 101 102 103 210 104 209 257 258 cell_2rw
* cell instance $1315 m0 *1 11.75,68.77
X$1315 101 102 103 218 104 220 257 258 cell_2rw
* cell instance $1316 r0 *1 11.75,65.78
X$1316 101 102 103 216 104 215 257 258 cell_2rw
* cell instance $1317 r0 *1 11.75,68.77
X$1317 101 102 103 224 104 223 257 258 cell_2rw
* cell instance $1318 m0 *1 11.75,71.76
X$1318 101 102 103 221 104 222 257 258 cell_2rw
* cell instance $1319 r0 *1 11.75,71.76
X$1319 101 102 103 226 104 225 257 258 cell_2rw
* cell instance $1320 m0 *1 11.75,74.75
X$1320 101 102 103 231 104 232 257 258 cell_2rw
* cell instance $1321 r0 *1 11.75,74.75
X$1321 101 102 103 230 104 229 257 258 cell_2rw
* cell instance $1322 m0 *1 11.75,77.74
X$1322 101 102 103 227 104 228 257 258 cell_2rw
* cell instance $1323 r0 *1 11.75,77.74
X$1323 101 102 103 237 104 238 257 258 cell_2rw
* cell instance $1324 m0 *1 11.75,80.73
X$1324 101 102 103 233 104 236 257 258 cell_2rw
* cell instance $1325 r0 *1 11.75,80.73
X$1325 101 102 103 235 104 234 257 258 cell_2rw
* cell instance $1326 m0 *1 11.75,83.72
X$1326 101 102 103 240 104 242 257 258 cell_2rw
* cell instance $1327 m0 *1 11.75,86.71
X$1327 101 102 103 244 104 243 257 258 cell_2rw
* cell instance $1328 r0 *1 11.75,83.72
X$1328 101 102 103 239 104 241 257 258 cell_2rw
* cell instance $1329 r0 *1 11.75,86.71
X$1329 101 102 103 245 104 247 257 258 cell_2rw
* cell instance $1330 m0 *1 11.75,89.7
X$1330 101 102 103 250 104 249 257 258 cell_2rw
* cell instance $1331 r0 *1 11.75,89.7
X$1331 101 102 103 246 104 248 257 258 cell_2rw
* cell instance $1332 m0 *1 11.75,92.69
X$1332 101 102 103 253 104 256 257 258 cell_2rw
* cell instance $1333 r0 *1 11.75,92.69
X$1333 101 102 103 255 104 254 257 258 cell_2rw
* cell instance $1334 m0 *1 11.75,95.68
X$1334 101 102 103 251 104 252 257 258 cell_2rw
* cell instance $1335 r0 *1 12.925,44.85
X$1335 105 106 107 127 108 128 257 258 cell_2rw
* cell instance $1336 m0 *1 12.925,47.84
X$1336 105 106 107 126 108 125 257 258 cell_2rw
* cell instance $1337 m0 *1 12.925,50.83
X$1337 105 106 107 195 108 197 257 258 cell_2rw
* cell instance $1338 r0 *1 12.925,47.84
X$1338 105 106 107 199 108 201 257 258 cell_2rw
* cell instance $1339 m0 *1 12.925,53.82
X$1339 105 106 107 198 108 193 257 258 cell_2rw
* cell instance $1340 r0 *1 12.925,50.83
X$1340 105 106 107 202 108 194 257 258 cell_2rw
* cell instance $1341 r0 *1 12.925,53.82
X$1341 105 106 107 196 108 200 257 258 cell_2rw
* cell instance $1342 m0 *1 12.925,56.81
X$1342 105 106 107 203 108 207 257 258 cell_2rw
* cell instance $1343 r0 *1 12.925,56.81
X$1343 105 106 107 206 108 208 257 258 cell_2rw
* cell instance $1344 m0 *1 12.925,59.8
X$1344 105 106 107 205 108 204 257 258 cell_2rw
* cell instance $1345 r0 *1 12.925,59.8
X$1345 105 106 107 214 108 213 257 258 cell_2rw
* cell instance $1346 m0 *1 12.925,62.79
X$1346 105 106 107 212 108 211 257 258 cell_2rw
* cell instance $1347 r0 *1 12.925,62.79
X$1347 105 106 107 210 108 209 257 258 cell_2rw
* cell instance $1348 m0 *1 12.925,65.78
X$1348 105 106 107 219 108 217 257 258 cell_2rw
* cell instance $1349 r0 *1 12.925,65.78
X$1349 105 106 107 216 108 215 257 258 cell_2rw
* cell instance $1350 m0 *1 12.925,68.77
X$1350 105 106 107 218 108 220 257 258 cell_2rw
* cell instance $1351 r0 *1 12.925,68.77
X$1351 105 106 107 224 108 223 257 258 cell_2rw
* cell instance $1352 m0 *1 12.925,71.76
X$1352 105 106 107 221 108 222 257 258 cell_2rw
* cell instance $1353 r0 *1 12.925,71.76
X$1353 105 106 107 226 108 225 257 258 cell_2rw
* cell instance $1354 m0 *1 12.925,74.75
X$1354 105 106 107 231 108 232 257 258 cell_2rw
* cell instance $1355 r0 *1 12.925,74.75
X$1355 105 106 107 230 108 229 257 258 cell_2rw
* cell instance $1356 m0 *1 12.925,77.74
X$1356 105 106 107 227 108 228 257 258 cell_2rw
* cell instance $1357 r0 *1 12.925,77.74
X$1357 105 106 107 237 108 238 257 258 cell_2rw
* cell instance $1358 m0 *1 12.925,80.73
X$1358 105 106 107 233 108 236 257 258 cell_2rw
* cell instance $1359 r0 *1 12.925,80.73
X$1359 105 106 107 235 108 234 257 258 cell_2rw
* cell instance $1360 m0 *1 12.925,83.72
X$1360 105 106 107 240 108 242 257 258 cell_2rw
* cell instance $1361 r0 *1 12.925,83.72
X$1361 105 106 107 239 108 241 257 258 cell_2rw
* cell instance $1362 m0 *1 12.925,86.71
X$1362 105 106 107 244 108 243 257 258 cell_2rw
* cell instance $1363 r0 *1 12.925,86.71
X$1363 105 106 107 245 108 247 257 258 cell_2rw
* cell instance $1364 m0 *1 12.925,89.7
X$1364 105 106 107 250 108 249 257 258 cell_2rw
* cell instance $1365 r0 *1 12.925,89.7
X$1365 105 106 107 246 108 248 257 258 cell_2rw
* cell instance $1366 m0 *1 12.925,92.69
X$1366 105 106 107 253 108 256 257 258 cell_2rw
* cell instance $1367 r0 *1 12.925,92.69
X$1367 105 106 107 255 108 254 257 258 cell_2rw
* cell instance $1368 m0 *1 12.925,95.68
X$1368 105 106 107 251 108 252 257 258 cell_2rw
* cell instance $1369 r0 *1 14.1,44.85
X$1369 109 110 111 127 112 128 257 258 cell_2rw
* cell instance $1370 m0 *1 14.1,47.84
X$1370 109 110 111 126 112 125 257 258 cell_2rw
* cell instance $1371 r0 *1 14.1,47.84
X$1371 109 110 111 199 112 201 257 258 cell_2rw
* cell instance $1372 m0 *1 14.1,50.83
X$1372 109 110 111 195 112 197 257 258 cell_2rw
* cell instance $1373 r0 *1 14.1,50.83
X$1373 109 110 111 202 112 194 257 258 cell_2rw
* cell instance $1374 m0 *1 14.1,53.82
X$1374 109 110 111 198 112 193 257 258 cell_2rw
* cell instance $1375 r0 *1 14.1,53.82
X$1375 109 110 111 196 112 200 257 258 cell_2rw
* cell instance $1376 m0 *1 14.1,56.81
X$1376 109 110 111 203 112 207 257 258 cell_2rw
* cell instance $1377 r0 *1 14.1,56.81
X$1377 109 110 111 206 112 208 257 258 cell_2rw
* cell instance $1378 m0 *1 14.1,59.8
X$1378 109 110 111 205 112 204 257 258 cell_2rw
* cell instance $1379 m0 *1 14.1,62.79
X$1379 109 110 111 212 112 211 257 258 cell_2rw
* cell instance $1380 r0 *1 14.1,59.8
X$1380 109 110 111 214 112 213 257 258 cell_2rw
* cell instance $1381 r0 *1 14.1,62.79
X$1381 109 110 111 210 112 209 257 258 cell_2rw
* cell instance $1382 m0 *1 14.1,65.78
X$1382 109 110 111 219 112 217 257 258 cell_2rw
* cell instance $1383 r0 *1 14.1,65.78
X$1383 109 110 111 216 112 215 257 258 cell_2rw
* cell instance $1384 m0 *1 14.1,68.77
X$1384 109 110 111 218 112 220 257 258 cell_2rw
* cell instance $1385 r0 *1 14.1,68.77
X$1385 109 110 111 224 112 223 257 258 cell_2rw
* cell instance $1386 m0 *1 14.1,71.76
X$1386 109 110 111 221 112 222 257 258 cell_2rw
* cell instance $1387 r0 *1 14.1,71.76
X$1387 109 110 111 226 112 225 257 258 cell_2rw
* cell instance $1388 m0 *1 14.1,74.75
X$1388 109 110 111 231 112 232 257 258 cell_2rw
* cell instance $1389 r0 *1 14.1,74.75
X$1389 109 110 111 230 112 229 257 258 cell_2rw
* cell instance $1390 m0 *1 14.1,77.74
X$1390 109 110 111 227 112 228 257 258 cell_2rw
* cell instance $1391 r0 *1 14.1,77.74
X$1391 109 110 111 237 112 238 257 258 cell_2rw
* cell instance $1392 m0 *1 14.1,80.73
X$1392 109 110 111 233 112 236 257 258 cell_2rw
* cell instance $1393 r0 *1 14.1,80.73
X$1393 109 110 111 235 112 234 257 258 cell_2rw
* cell instance $1394 m0 *1 14.1,83.72
X$1394 109 110 111 240 112 242 257 258 cell_2rw
* cell instance $1395 m0 *1 14.1,86.71
X$1395 109 110 111 244 112 243 257 258 cell_2rw
* cell instance $1396 r0 *1 14.1,83.72
X$1396 109 110 111 239 112 241 257 258 cell_2rw
* cell instance $1397 r0 *1 14.1,86.71
X$1397 109 110 111 245 112 247 257 258 cell_2rw
* cell instance $1398 m0 *1 14.1,89.7
X$1398 109 110 111 250 112 249 257 258 cell_2rw
* cell instance $1399 r0 *1 14.1,89.7
X$1399 109 110 111 246 112 248 257 258 cell_2rw
* cell instance $1400 m0 *1 14.1,92.69
X$1400 109 110 111 253 112 256 257 258 cell_2rw
* cell instance $1401 r0 *1 14.1,92.69
X$1401 109 110 111 255 112 254 257 258 cell_2rw
* cell instance $1402 m0 *1 14.1,95.68
X$1402 109 110 111 251 112 252 257 258 cell_2rw
* cell instance $1403 r0 *1 15.275,44.85
X$1403 113 114 115 127 116 128 257 258 cell_2rw
* cell instance $1404 m0 *1 15.275,47.84
X$1404 113 114 115 126 116 125 257 258 cell_2rw
* cell instance $1405 m0 *1 15.275,50.83
X$1405 113 114 115 195 116 197 257 258 cell_2rw
* cell instance $1406 r0 *1 15.275,47.84
X$1406 113 114 115 199 116 201 257 258 cell_2rw
* cell instance $1407 m0 *1 15.275,53.82
X$1407 113 114 115 198 116 193 257 258 cell_2rw
* cell instance $1408 r0 *1 15.275,50.83
X$1408 113 114 115 202 116 194 257 258 cell_2rw
* cell instance $1409 r0 *1 15.275,53.82
X$1409 113 114 115 196 116 200 257 258 cell_2rw
* cell instance $1410 m0 *1 15.275,56.81
X$1410 113 114 115 203 116 207 257 258 cell_2rw
* cell instance $1411 r0 *1 15.275,56.81
X$1411 113 114 115 206 116 208 257 258 cell_2rw
* cell instance $1412 m0 *1 15.275,59.8
X$1412 113 114 115 205 116 204 257 258 cell_2rw
* cell instance $1413 r0 *1 15.275,59.8
X$1413 113 114 115 214 116 213 257 258 cell_2rw
* cell instance $1414 m0 *1 15.275,62.79
X$1414 113 114 115 212 116 211 257 258 cell_2rw
* cell instance $1415 r0 *1 15.275,62.79
X$1415 113 114 115 210 116 209 257 258 cell_2rw
* cell instance $1416 m0 *1 15.275,65.78
X$1416 113 114 115 219 116 217 257 258 cell_2rw
* cell instance $1417 r0 *1 15.275,65.78
X$1417 113 114 115 216 116 215 257 258 cell_2rw
* cell instance $1418 m0 *1 15.275,68.77
X$1418 113 114 115 218 116 220 257 258 cell_2rw
* cell instance $1419 r0 *1 15.275,68.77
X$1419 113 114 115 224 116 223 257 258 cell_2rw
* cell instance $1420 m0 *1 15.275,71.76
X$1420 113 114 115 221 116 222 257 258 cell_2rw
* cell instance $1421 r0 *1 15.275,71.76
X$1421 113 114 115 226 116 225 257 258 cell_2rw
* cell instance $1422 m0 *1 15.275,74.75
X$1422 113 114 115 231 116 232 257 258 cell_2rw
* cell instance $1423 r0 *1 15.275,74.75
X$1423 113 114 115 230 116 229 257 258 cell_2rw
* cell instance $1424 m0 *1 15.275,77.74
X$1424 113 114 115 227 116 228 257 258 cell_2rw
* cell instance $1425 m0 *1 15.275,80.73
X$1425 113 114 115 233 116 236 257 258 cell_2rw
* cell instance $1426 r0 *1 15.275,77.74
X$1426 113 114 115 237 116 238 257 258 cell_2rw
* cell instance $1427 m0 *1 15.275,83.72
X$1427 113 114 115 240 116 242 257 258 cell_2rw
* cell instance $1428 r0 *1 15.275,80.73
X$1428 113 114 115 235 116 234 257 258 cell_2rw
* cell instance $1429 r0 *1 15.275,83.72
X$1429 113 114 115 239 116 241 257 258 cell_2rw
* cell instance $1430 m0 *1 15.275,86.71
X$1430 113 114 115 244 116 243 257 258 cell_2rw
* cell instance $1431 m0 *1 15.275,89.7
X$1431 113 114 115 250 116 249 257 258 cell_2rw
* cell instance $1432 r0 *1 15.275,86.71
X$1432 113 114 115 245 116 247 257 258 cell_2rw
* cell instance $1433 r0 *1 15.275,89.7
X$1433 113 114 115 246 116 248 257 258 cell_2rw
* cell instance $1434 m0 *1 15.275,92.69
X$1434 113 114 115 253 116 256 257 258 cell_2rw
* cell instance $1435 r0 *1 15.275,92.69
X$1435 113 114 115 255 116 254 257 258 cell_2rw
* cell instance $1436 m0 *1 15.275,95.68
X$1436 113 114 115 251 116 252 257 258 cell_2rw
* cell instance $1437 r0 *1 16.45,44.85
X$1437 117 118 119 127 120 128 257 258 cell_2rw
* cell instance $1438 m0 *1 16.45,47.84
X$1438 117 118 119 126 120 125 257 258 cell_2rw
* cell instance $1439 r0 *1 16.45,47.84
X$1439 117 118 119 199 120 201 257 258 cell_2rw
* cell instance $1440 m0 *1 16.45,50.83
X$1440 117 118 119 195 120 197 257 258 cell_2rw
* cell instance $1441 m0 *1 16.45,53.82
X$1441 117 118 119 198 120 193 257 258 cell_2rw
* cell instance $1442 r0 *1 16.45,50.83
X$1442 117 118 119 202 120 194 257 258 cell_2rw
* cell instance $1443 r0 *1 16.45,53.82
X$1443 117 118 119 196 120 200 257 258 cell_2rw
* cell instance $1444 m0 *1 16.45,56.81
X$1444 117 118 119 203 120 207 257 258 cell_2rw
* cell instance $1445 m0 *1 16.45,59.8
X$1445 117 118 119 205 120 204 257 258 cell_2rw
* cell instance $1446 r0 *1 16.45,56.81
X$1446 117 118 119 206 120 208 257 258 cell_2rw
* cell instance $1447 m0 *1 16.45,62.79
X$1447 117 118 119 212 120 211 257 258 cell_2rw
* cell instance $1448 r0 *1 16.45,59.8
X$1448 117 118 119 214 120 213 257 258 cell_2rw
* cell instance $1449 r0 *1 16.45,62.79
X$1449 117 118 119 210 120 209 257 258 cell_2rw
* cell instance $1450 m0 *1 16.45,65.78
X$1450 117 118 119 219 120 217 257 258 cell_2rw
* cell instance $1451 r0 *1 16.45,65.78
X$1451 117 118 119 216 120 215 257 258 cell_2rw
* cell instance $1452 m0 *1 16.45,68.77
X$1452 117 118 119 218 120 220 257 258 cell_2rw
* cell instance $1453 r0 *1 16.45,68.77
X$1453 117 118 119 224 120 223 257 258 cell_2rw
* cell instance $1454 m0 *1 16.45,71.76
X$1454 117 118 119 221 120 222 257 258 cell_2rw
* cell instance $1455 r0 *1 16.45,71.76
X$1455 117 118 119 226 120 225 257 258 cell_2rw
* cell instance $1456 m0 *1 16.45,74.75
X$1456 117 118 119 231 120 232 257 258 cell_2rw
* cell instance $1457 r0 *1 16.45,74.75
X$1457 117 118 119 230 120 229 257 258 cell_2rw
* cell instance $1458 m0 *1 16.45,77.74
X$1458 117 118 119 227 120 228 257 258 cell_2rw
* cell instance $1459 m0 *1 16.45,80.73
X$1459 117 118 119 233 120 236 257 258 cell_2rw
* cell instance $1460 r0 *1 16.45,77.74
X$1460 117 118 119 237 120 238 257 258 cell_2rw
* cell instance $1461 r0 *1 16.45,80.73
X$1461 117 118 119 235 120 234 257 258 cell_2rw
* cell instance $1462 m0 *1 16.45,83.72
X$1462 117 118 119 240 120 242 257 258 cell_2rw
* cell instance $1463 r0 *1 16.45,83.72
X$1463 117 118 119 239 120 241 257 258 cell_2rw
* cell instance $1464 m0 *1 16.45,86.71
X$1464 117 118 119 244 120 243 257 258 cell_2rw
* cell instance $1465 r0 *1 16.45,86.71
X$1465 117 118 119 245 120 247 257 258 cell_2rw
* cell instance $1466 m0 *1 16.45,89.7
X$1466 117 118 119 250 120 249 257 258 cell_2rw
* cell instance $1467 r0 *1 16.45,89.7
X$1467 117 118 119 246 120 248 257 258 cell_2rw
* cell instance $1468 m0 *1 16.45,92.69
X$1468 117 118 119 253 120 256 257 258 cell_2rw
* cell instance $1469 r0 *1 16.45,92.69
X$1469 117 118 119 255 120 254 257 258 cell_2rw
* cell instance $1470 m0 *1 16.45,95.68
X$1470 117 118 119 251 120 252 257 258 cell_2rw
* cell instance $1471 r0 *1 17.625,44.85
X$1471 121 122 123 127 124 128 257 258 cell_2rw
* cell instance $1472 m0 *1 17.625,47.84
X$1472 121 122 123 126 124 125 257 258 cell_2rw
* cell instance $1473 m0 *1 17.625,50.83
X$1473 121 122 123 195 124 197 257 258 cell_2rw
* cell instance $1474 r0 *1 17.625,47.84
X$1474 121 122 123 199 124 201 257 258 cell_2rw
* cell instance $1475 r0 *1 17.625,50.83
X$1475 121 122 123 202 124 194 257 258 cell_2rw
* cell instance $1476 m0 *1 17.625,53.82
X$1476 121 122 123 198 124 193 257 258 cell_2rw
* cell instance $1477 m0 *1 17.625,56.81
X$1477 121 122 123 203 124 207 257 258 cell_2rw
* cell instance $1478 r0 *1 17.625,53.82
X$1478 121 122 123 196 124 200 257 258 cell_2rw
* cell instance $1479 m0 *1 17.625,59.8
X$1479 121 122 123 205 124 204 257 258 cell_2rw
* cell instance $1480 r0 *1 17.625,56.81
X$1480 121 122 123 206 124 208 257 258 cell_2rw
* cell instance $1481 m0 *1 17.625,62.79
X$1481 121 122 123 212 124 211 257 258 cell_2rw
* cell instance $1482 r0 *1 17.625,59.8
X$1482 121 122 123 214 124 213 257 258 cell_2rw
* cell instance $1483 m0 *1 17.625,65.78
X$1483 121 122 123 219 124 217 257 258 cell_2rw
* cell instance $1484 r0 *1 17.625,62.79
X$1484 121 122 123 210 124 209 257 258 cell_2rw
* cell instance $1485 r0 *1 17.625,65.78
X$1485 121 122 123 216 124 215 257 258 cell_2rw
* cell instance $1486 m0 *1 17.625,68.77
X$1486 121 122 123 218 124 220 257 258 cell_2rw
* cell instance $1487 m0 *1 17.625,71.76
X$1487 121 122 123 221 124 222 257 258 cell_2rw
* cell instance $1488 r0 *1 17.625,68.77
X$1488 121 122 123 224 124 223 257 258 cell_2rw
* cell instance $1489 r0 *1 17.625,71.76
X$1489 121 122 123 226 124 225 257 258 cell_2rw
* cell instance $1490 m0 *1 17.625,74.75
X$1490 121 122 123 231 124 232 257 258 cell_2rw
* cell instance $1491 r0 *1 17.625,74.75
X$1491 121 122 123 230 124 229 257 258 cell_2rw
* cell instance $1492 m0 *1 17.625,77.74
X$1492 121 122 123 227 124 228 257 258 cell_2rw
* cell instance $1493 r0 *1 17.625,77.74
X$1493 121 122 123 237 124 238 257 258 cell_2rw
* cell instance $1494 m0 *1 17.625,80.73
X$1494 121 122 123 233 124 236 257 258 cell_2rw
* cell instance $1495 r0 *1 17.625,80.73
X$1495 121 122 123 235 124 234 257 258 cell_2rw
* cell instance $1496 m0 *1 17.625,83.72
X$1496 121 122 123 240 124 242 257 258 cell_2rw
* cell instance $1497 r0 *1 17.625,83.72
X$1497 121 122 123 239 124 241 257 258 cell_2rw
* cell instance $1498 m0 *1 17.625,86.71
X$1498 121 122 123 244 124 243 257 258 cell_2rw
* cell instance $1499 r0 *1 17.625,86.71
X$1499 121 122 123 245 124 247 257 258 cell_2rw
* cell instance $1500 m0 *1 17.625,89.7
X$1500 121 122 123 250 124 249 257 258 cell_2rw
* cell instance $1501 m0 *1 17.625,92.69
X$1501 121 122 123 253 124 256 257 258 cell_2rw
* cell instance $1502 r0 *1 17.625,89.7
X$1502 121 122 123 246 124 248 257 258 cell_2rw
* cell instance $1503 m0 *1 17.625,95.68
X$1503 121 122 123 251 124 252 257 258 cell_2rw
* cell instance $1504 r0 *1 17.625,92.69
X$1504 121 122 123 255 124 254 257 258 cell_2rw
* cell instance $1505 m0 *1 18.8,47.84
X$1505 129 130 131 126 132 125 257 258 cell_2rw
* cell instance $1506 m0 *1 19.975,47.84
X$1506 133 134 135 126 136 125 257 258 cell_2rw
* cell instance $1507 m0 *1 21.15,47.84
X$1507 137 138 139 126 140 125 257 258 cell_2rw
* cell instance $1508 m0 *1 22.325,47.84
X$1508 141 142 143 126 144 125 257 258 cell_2rw
* cell instance $1509 m0 *1 23.5,47.84
X$1509 145 146 147 126 148 125 257 258 cell_2rw
* cell instance $1510 m0 *1 24.675,47.84
X$1510 149 150 151 126 152 125 257 258 cell_2rw
* cell instance $1511 m0 *1 25.85,47.84
X$1511 153 154 155 126 156 125 257 258 cell_2rw
* cell instance $1512 m0 *1 27.025,47.84
X$1512 157 158 159 126 160 125 257 258 cell_2rw
* cell instance $1513 m0 *1 28.2,47.84
X$1513 161 162 163 126 164 125 257 258 cell_2rw
* cell instance $1514 m0 *1 29.375,47.84
X$1514 165 166 167 126 168 125 257 258 cell_2rw
* cell instance $1515 m0 *1 30.55,47.84
X$1515 169 170 171 126 172 125 257 258 cell_2rw
* cell instance $1516 m0 *1 31.725,47.84
X$1516 173 174 175 126 176 125 257 258 cell_2rw
* cell instance $1517 m0 *1 32.9,47.84
X$1517 177 178 179 126 180 125 257 258 cell_2rw
* cell instance $1518 m0 *1 34.075,47.84
X$1518 181 182 183 126 184 125 257 258 cell_2rw
* cell instance $1519 m0 *1 35.25,47.84
X$1519 185 186 187 126 188 125 257 258 cell_2rw
* cell instance $1520 m0 *1 36.425,47.84
X$1520 189 190 191 126 192 125 257 258 cell_2rw
* cell instance $1521 r0 *1 18.8,44.85
X$1521 129 130 131 127 132 128 257 258 cell_2rw
* cell instance $1522 r0 *1 19.975,44.85
X$1522 133 134 135 127 136 128 257 258 cell_2rw
* cell instance $1523 r0 *1 21.15,44.85
X$1523 137 138 139 127 140 128 257 258 cell_2rw
* cell instance $1524 r0 *1 22.325,44.85
X$1524 141 142 143 127 144 128 257 258 cell_2rw
* cell instance $1525 r0 *1 23.5,44.85
X$1525 145 146 147 127 148 128 257 258 cell_2rw
* cell instance $1526 r0 *1 24.675,44.85
X$1526 149 150 151 127 152 128 257 258 cell_2rw
* cell instance $1527 r0 *1 25.85,44.85
X$1527 153 154 155 127 156 128 257 258 cell_2rw
* cell instance $1528 r0 *1 27.025,44.85
X$1528 157 158 159 127 160 128 257 258 cell_2rw
* cell instance $1529 r0 *1 28.2,44.85
X$1529 161 162 163 127 164 128 257 258 cell_2rw
* cell instance $1530 r0 *1 29.375,44.85
X$1530 165 166 167 127 168 128 257 258 cell_2rw
* cell instance $1531 r0 *1 30.55,44.85
X$1531 169 170 171 127 172 128 257 258 cell_2rw
* cell instance $1532 r0 *1 31.725,44.85
X$1532 173 174 175 127 176 128 257 258 cell_2rw
* cell instance $1533 r0 *1 32.9,44.85
X$1533 177 178 179 127 180 128 257 258 cell_2rw
* cell instance $1534 r0 *1 34.075,44.85
X$1534 181 182 183 127 184 128 257 258 cell_2rw
* cell instance $1535 r0 *1 35.25,44.85
X$1535 185 186 187 127 188 128 257 258 cell_2rw
* cell instance $1536 r0 *1 36.425,44.85
X$1536 189 190 191 127 192 128 257 258 cell_2rw
* cell instance $1537 r0 *1 18.8,47.84
X$1537 129 130 131 199 132 201 257 258 cell_2rw
* cell instance $1538 m0 *1 18.8,50.83
X$1538 129 130 131 195 132 197 257 258 cell_2rw
* cell instance $1539 r0 *1 18.8,50.83
X$1539 129 130 131 202 132 194 257 258 cell_2rw
* cell instance $1540 m0 *1 18.8,53.82
X$1540 129 130 131 198 132 193 257 258 cell_2rw
* cell instance $1541 r0 *1 18.8,53.82
X$1541 129 130 131 196 132 200 257 258 cell_2rw
* cell instance $1542 m0 *1 18.8,56.81
X$1542 129 130 131 203 132 207 257 258 cell_2rw
* cell instance $1543 r0 *1 18.8,56.81
X$1543 129 130 131 206 132 208 257 258 cell_2rw
* cell instance $1544 m0 *1 18.8,59.8
X$1544 129 130 131 205 132 204 257 258 cell_2rw
* cell instance $1545 r0 *1 18.8,59.8
X$1545 129 130 131 214 132 213 257 258 cell_2rw
* cell instance $1546 m0 *1 18.8,62.79
X$1546 129 130 131 212 132 211 257 258 cell_2rw
* cell instance $1547 r0 *1 18.8,62.79
X$1547 129 130 131 210 132 209 257 258 cell_2rw
* cell instance $1548 m0 *1 18.8,65.78
X$1548 129 130 131 219 132 217 257 258 cell_2rw
* cell instance $1549 r0 *1 18.8,65.78
X$1549 129 130 131 216 132 215 257 258 cell_2rw
* cell instance $1550 m0 *1 18.8,68.77
X$1550 129 130 131 218 132 220 257 258 cell_2rw
* cell instance $1551 m0 *1 18.8,71.76
X$1551 129 130 131 221 132 222 257 258 cell_2rw
* cell instance $1552 r0 *1 18.8,68.77
X$1552 129 130 131 224 132 223 257 258 cell_2rw
* cell instance $1553 m0 *1 18.8,74.75
X$1553 129 130 131 231 132 232 257 258 cell_2rw
* cell instance $1554 r0 *1 18.8,71.76
X$1554 129 130 131 226 132 225 257 258 cell_2rw
* cell instance $1555 m0 *1 18.8,77.74
X$1555 129 130 131 227 132 228 257 258 cell_2rw
* cell instance $1556 r0 *1 18.8,74.75
X$1556 129 130 131 230 132 229 257 258 cell_2rw
* cell instance $1557 r0 *1 18.8,77.74
X$1557 129 130 131 237 132 238 257 258 cell_2rw
* cell instance $1558 m0 *1 18.8,80.73
X$1558 129 130 131 233 132 236 257 258 cell_2rw
* cell instance $1559 r0 *1 18.8,80.73
X$1559 129 130 131 235 132 234 257 258 cell_2rw
* cell instance $1560 m0 *1 18.8,83.72
X$1560 129 130 131 240 132 242 257 258 cell_2rw
* cell instance $1561 r0 *1 18.8,83.72
X$1561 129 130 131 239 132 241 257 258 cell_2rw
* cell instance $1562 m0 *1 18.8,86.71
X$1562 129 130 131 244 132 243 257 258 cell_2rw
* cell instance $1563 r0 *1 18.8,86.71
X$1563 129 130 131 245 132 247 257 258 cell_2rw
* cell instance $1564 m0 *1 18.8,89.7
X$1564 129 130 131 250 132 249 257 258 cell_2rw
* cell instance $1565 r0 *1 18.8,89.7
X$1565 129 130 131 246 132 248 257 258 cell_2rw
* cell instance $1566 m0 *1 18.8,92.69
X$1566 129 130 131 253 132 256 257 258 cell_2rw
* cell instance $1567 r0 *1 18.8,92.69
X$1567 129 130 131 255 132 254 257 258 cell_2rw
* cell instance $1568 m0 *1 18.8,95.68
X$1568 129 130 131 251 132 252 257 258 cell_2rw
* cell instance $1569 r0 *1 19.975,47.84
X$1569 133 134 135 199 136 201 257 258 cell_2rw
* cell instance $1570 m0 *1 19.975,50.83
X$1570 133 134 135 195 136 197 257 258 cell_2rw
* cell instance $1571 r0 *1 19.975,50.83
X$1571 133 134 135 202 136 194 257 258 cell_2rw
* cell instance $1572 m0 *1 19.975,53.82
X$1572 133 134 135 198 136 193 257 258 cell_2rw
* cell instance $1573 m0 *1 19.975,56.81
X$1573 133 134 135 203 136 207 257 258 cell_2rw
* cell instance $1574 r0 *1 19.975,53.82
X$1574 133 134 135 196 136 200 257 258 cell_2rw
* cell instance $1575 r0 *1 19.975,56.81
X$1575 133 134 135 206 136 208 257 258 cell_2rw
* cell instance $1576 m0 *1 19.975,59.8
X$1576 133 134 135 205 136 204 257 258 cell_2rw
* cell instance $1577 r0 *1 19.975,59.8
X$1577 133 134 135 214 136 213 257 258 cell_2rw
* cell instance $1578 m0 *1 19.975,62.79
X$1578 133 134 135 212 136 211 257 258 cell_2rw
* cell instance $1579 r0 *1 19.975,62.79
X$1579 133 134 135 210 136 209 257 258 cell_2rw
* cell instance $1580 m0 *1 19.975,65.78
X$1580 133 134 135 219 136 217 257 258 cell_2rw
* cell instance $1581 r0 *1 19.975,65.78
X$1581 133 134 135 216 136 215 257 258 cell_2rw
* cell instance $1582 m0 *1 19.975,68.77
X$1582 133 134 135 218 136 220 257 258 cell_2rw
* cell instance $1583 r0 *1 19.975,68.77
X$1583 133 134 135 224 136 223 257 258 cell_2rw
* cell instance $1584 m0 *1 19.975,71.76
X$1584 133 134 135 221 136 222 257 258 cell_2rw
* cell instance $1585 r0 *1 19.975,71.76
X$1585 133 134 135 226 136 225 257 258 cell_2rw
* cell instance $1586 m0 *1 19.975,74.75
X$1586 133 134 135 231 136 232 257 258 cell_2rw
* cell instance $1587 r0 *1 19.975,74.75
X$1587 133 134 135 230 136 229 257 258 cell_2rw
* cell instance $1588 m0 *1 19.975,77.74
X$1588 133 134 135 227 136 228 257 258 cell_2rw
* cell instance $1589 m0 *1 19.975,80.73
X$1589 133 134 135 233 136 236 257 258 cell_2rw
* cell instance $1590 r0 *1 19.975,77.74
X$1590 133 134 135 237 136 238 257 258 cell_2rw
* cell instance $1591 r0 *1 19.975,80.73
X$1591 133 134 135 235 136 234 257 258 cell_2rw
* cell instance $1592 m0 *1 19.975,83.72
X$1592 133 134 135 240 136 242 257 258 cell_2rw
* cell instance $1593 r0 *1 19.975,83.72
X$1593 133 134 135 239 136 241 257 258 cell_2rw
* cell instance $1594 m0 *1 19.975,86.71
X$1594 133 134 135 244 136 243 257 258 cell_2rw
* cell instance $1595 r0 *1 19.975,86.71
X$1595 133 134 135 245 136 247 257 258 cell_2rw
* cell instance $1596 m0 *1 19.975,89.7
X$1596 133 134 135 250 136 249 257 258 cell_2rw
* cell instance $1597 r0 *1 19.975,89.7
X$1597 133 134 135 246 136 248 257 258 cell_2rw
* cell instance $1598 m0 *1 19.975,92.69
X$1598 133 134 135 253 136 256 257 258 cell_2rw
* cell instance $1599 r0 *1 19.975,92.69
X$1599 133 134 135 255 136 254 257 258 cell_2rw
* cell instance $1600 m0 *1 19.975,95.68
X$1600 133 134 135 251 136 252 257 258 cell_2rw
* cell instance $1601 r0 *1 21.15,47.84
X$1601 137 138 139 199 140 201 257 258 cell_2rw
* cell instance $1602 m0 *1 21.15,50.83
X$1602 137 138 139 195 140 197 257 258 cell_2rw
* cell instance $1603 r0 *1 21.15,50.83
X$1603 137 138 139 202 140 194 257 258 cell_2rw
* cell instance $1604 m0 *1 21.15,53.82
X$1604 137 138 139 198 140 193 257 258 cell_2rw
* cell instance $1605 r0 *1 21.15,53.82
X$1605 137 138 139 196 140 200 257 258 cell_2rw
* cell instance $1606 m0 *1 21.15,56.81
X$1606 137 138 139 203 140 207 257 258 cell_2rw
* cell instance $1607 r0 *1 21.15,56.81
X$1607 137 138 139 206 140 208 257 258 cell_2rw
* cell instance $1608 m0 *1 21.15,59.8
X$1608 137 138 139 205 140 204 257 258 cell_2rw
* cell instance $1609 r0 *1 21.15,59.8
X$1609 137 138 139 214 140 213 257 258 cell_2rw
* cell instance $1610 m0 *1 21.15,62.79
X$1610 137 138 139 212 140 211 257 258 cell_2rw
* cell instance $1611 r0 *1 21.15,62.79
X$1611 137 138 139 210 140 209 257 258 cell_2rw
* cell instance $1612 m0 *1 21.15,65.78
X$1612 137 138 139 219 140 217 257 258 cell_2rw
* cell instance $1613 r0 *1 21.15,65.78
X$1613 137 138 139 216 140 215 257 258 cell_2rw
* cell instance $1614 m0 *1 21.15,68.77
X$1614 137 138 139 218 140 220 257 258 cell_2rw
* cell instance $1615 r0 *1 21.15,68.77
X$1615 137 138 139 224 140 223 257 258 cell_2rw
* cell instance $1616 m0 *1 21.15,71.76
X$1616 137 138 139 221 140 222 257 258 cell_2rw
* cell instance $1617 r0 *1 21.15,71.76
X$1617 137 138 139 226 140 225 257 258 cell_2rw
* cell instance $1618 m0 *1 21.15,74.75
X$1618 137 138 139 231 140 232 257 258 cell_2rw
* cell instance $1619 r0 *1 21.15,74.75
X$1619 137 138 139 230 140 229 257 258 cell_2rw
* cell instance $1620 m0 *1 21.15,77.74
X$1620 137 138 139 227 140 228 257 258 cell_2rw
* cell instance $1621 r0 *1 21.15,77.74
X$1621 137 138 139 237 140 238 257 258 cell_2rw
* cell instance $1622 m0 *1 21.15,80.73
X$1622 137 138 139 233 140 236 257 258 cell_2rw
* cell instance $1623 r0 *1 21.15,80.73
X$1623 137 138 139 235 140 234 257 258 cell_2rw
* cell instance $1624 m0 *1 21.15,83.72
X$1624 137 138 139 240 140 242 257 258 cell_2rw
* cell instance $1625 r0 *1 21.15,83.72
X$1625 137 138 139 239 140 241 257 258 cell_2rw
* cell instance $1626 m0 *1 21.15,86.71
X$1626 137 138 139 244 140 243 257 258 cell_2rw
* cell instance $1627 r0 *1 21.15,86.71
X$1627 137 138 139 245 140 247 257 258 cell_2rw
* cell instance $1628 m0 *1 21.15,89.7
X$1628 137 138 139 250 140 249 257 258 cell_2rw
* cell instance $1629 r0 *1 21.15,89.7
X$1629 137 138 139 246 140 248 257 258 cell_2rw
* cell instance $1630 m0 *1 21.15,92.69
X$1630 137 138 139 253 140 256 257 258 cell_2rw
* cell instance $1631 r0 *1 21.15,92.69
X$1631 137 138 139 255 140 254 257 258 cell_2rw
* cell instance $1632 m0 *1 21.15,95.68
X$1632 137 138 139 251 140 252 257 258 cell_2rw
* cell instance $1633 r0 *1 22.325,47.84
X$1633 141 142 143 199 144 201 257 258 cell_2rw
* cell instance $1634 m0 *1 22.325,50.83
X$1634 141 142 143 195 144 197 257 258 cell_2rw
* cell instance $1635 r0 *1 22.325,50.83
X$1635 141 142 143 202 144 194 257 258 cell_2rw
* cell instance $1636 m0 *1 22.325,53.82
X$1636 141 142 143 198 144 193 257 258 cell_2rw
* cell instance $1637 m0 *1 22.325,56.81
X$1637 141 142 143 203 144 207 257 258 cell_2rw
* cell instance $1638 r0 *1 22.325,53.82
X$1638 141 142 143 196 144 200 257 258 cell_2rw
* cell instance $1639 r0 *1 22.325,56.81
X$1639 141 142 143 206 144 208 257 258 cell_2rw
* cell instance $1640 m0 *1 22.325,59.8
X$1640 141 142 143 205 144 204 257 258 cell_2rw
* cell instance $1641 r0 *1 22.325,59.8
X$1641 141 142 143 214 144 213 257 258 cell_2rw
* cell instance $1642 m0 *1 22.325,62.79
X$1642 141 142 143 212 144 211 257 258 cell_2rw
* cell instance $1643 r0 *1 22.325,62.79
X$1643 141 142 143 210 144 209 257 258 cell_2rw
* cell instance $1644 m0 *1 22.325,65.78
X$1644 141 142 143 219 144 217 257 258 cell_2rw
* cell instance $1645 r0 *1 22.325,65.78
X$1645 141 142 143 216 144 215 257 258 cell_2rw
* cell instance $1646 m0 *1 22.325,68.77
X$1646 141 142 143 218 144 220 257 258 cell_2rw
* cell instance $1647 r0 *1 22.325,68.77
X$1647 141 142 143 224 144 223 257 258 cell_2rw
* cell instance $1648 m0 *1 22.325,71.76
X$1648 141 142 143 221 144 222 257 258 cell_2rw
* cell instance $1649 r0 *1 22.325,71.76
X$1649 141 142 143 226 144 225 257 258 cell_2rw
* cell instance $1650 m0 *1 22.325,74.75
X$1650 141 142 143 231 144 232 257 258 cell_2rw
* cell instance $1651 r0 *1 22.325,74.75
X$1651 141 142 143 230 144 229 257 258 cell_2rw
* cell instance $1652 m0 *1 22.325,77.74
X$1652 141 142 143 227 144 228 257 258 cell_2rw
* cell instance $1653 r0 *1 22.325,77.74
X$1653 141 142 143 237 144 238 257 258 cell_2rw
* cell instance $1654 m0 *1 22.325,80.73
X$1654 141 142 143 233 144 236 257 258 cell_2rw
* cell instance $1655 r0 *1 22.325,80.73
X$1655 141 142 143 235 144 234 257 258 cell_2rw
* cell instance $1656 m0 *1 22.325,83.72
X$1656 141 142 143 240 144 242 257 258 cell_2rw
* cell instance $1657 r0 *1 22.325,83.72
X$1657 141 142 143 239 144 241 257 258 cell_2rw
* cell instance $1658 m0 *1 22.325,86.71
X$1658 141 142 143 244 144 243 257 258 cell_2rw
* cell instance $1659 m0 *1 22.325,89.7
X$1659 141 142 143 250 144 249 257 258 cell_2rw
* cell instance $1660 r0 *1 22.325,86.71
X$1660 141 142 143 245 144 247 257 258 cell_2rw
* cell instance $1661 m0 *1 22.325,92.69
X$1661 141 142 143 253 144 256 257 258 cell_2rw
* cell instance $1662 r0 *1 22.325,89.7
X$1662 141 142 143 246 144 248 257 258 cell_2rw
* cell instance $1663 r0 *1 22.325,92.69
X$1663 141 142 143 255 144 254 257 258 cell_2rw
* cell instance $1664 m0 *1 22.325,95.68
X$1664 141 142 143 251 144 252 257 258 cell_2rw
* cell instance $1665 r0 *1 23.5,47.84
X$1665 145 146 147 199 148 201 257 258 cell_2rw
* cell instance $1666 m0 *1 23.5,50.83
X$1666 145 146 147 195 148 197 257 258 cell_2rw
* cell instance $1667 r0 *1 23.5,50.83
X$1667 145 146 147 202 148 194 257 258 cell_2rw
* cell instance $1668 m0 *1 23.5,53.82
X$1668 145 146 147 198 148 193 257 258 cell_2rw
* cell instance $1669 r0 *1 23.5,53.82
X$1669 145 146 147 196 148 200 257 258 cell_2rw
* cell instance $1670 m0 *1 23.5,56.81
X$1670 145 146 147 203 148 207 257 258 cell_2rw
* cell instance $1671 r0 *1 23.5,56.81
X$1671 145 146 147 206 148 208 257 258 cell_2rw
* cell instance $1672 m0 *1 23.5,59.8
X$1672 145 146 147 205 148 204 257 258 cell_2rw
* cell instance $1673 r0 *1 23.5,59.8
X$1673 145 146 147 214 148 213 257 258 cell_2rw
* cell instance $1674 m0 *1 23.5,62.79
X$1674 145 146 147 212 148 211 257 258 cell_2rw
* cell instance $1675 r0 *1 23.5,62.79
X$1675 145 146 147 210 148 209 257 258 cell_2rw
* cell instance $1676 m0 *1 23.5,65.78
X$1676 145 146 147 219 148 217 257 258 cell_2rw
* cell instance $1677 r0 *1 23.5,65.78
X$1677 145 146 147 216 148 215 257 258 cell_2rw
* cell instance $1678 m0 *1 23.5,68.77
X$1678 145 146 147 218 148 220 257 258 cell_2rw
* cell instance $1679 m0 *1 23.5,71.76
X$1679 145 146 147 221 148 222 257 258 cell_2rw
* cell instance $1680 r0 *1 23.5,68.77
X$1680 145 146 147 224 148 223 257 258 cell_2rw
* cell instance $1681 r0 *1 23.5,71.76
X$1681 145 146 147 226 148 225 257 258 cell_2rw
* cell instance $1682 m0 *1 23.5,74.75
X$1682 145 146 147 231 148 232 257 258 cell_2rw
* cell instance $1683 r0 *1 23.5,74.75
X$1683 145 146 147 230 148 229 257 258 cell_2rw
* cell instance $1684 m0 *1 23.5,77.74
X$1684 145 146 147 227 148 228 257 258 cell_2rw
* cell instance $1685 r0 *1 23.5,77.74
X$1685 145 146 147 237 148 238 257 258 cell_2rw
* cell instance $1686 m0 *1 23.5,80.73
X$1686 145 146 147 233 148 236 257 258 cell_2rw
* cell instance $1687 m0 *1 23.5,83.72
X$1687 145 146 147 240 148 242 257 258 cell_2rw
* cell instance $1688 r0 *1 23.5,80.73
X$1688 145 146 147 235 148 234 257 258 cell_2rw
* cell instance $1689 r0 *1 23.5,83.72
X$1689 145 146 147 239 148 241 257 258 cell_2rw
* cell instance $1690 m0 *1 23.5,86.71
X$1690 145 146 147 244 148 243 257 258 cell_2rw
* cell instance $1691 r0 *1 23.5,86.71
X$1691 145 146 147 245 148 247 257 258 cell_2rw
* cell instance $1692 m0 *1 23.5,89.7
X$1692 145 146 147 250 148 249 257 258 cell_2rw
* cell instance $1693 r0 *1 23.5,89.7
X$1693 145 146 147 246 148 248 257 258 cell_2rw
* cell instance $1694 m0 *1 23.5,92.69
X$1694 145 146 147 253 148 256 257 258 cell_2rw
* cell instance $1695 m0 *1 23.5,95.68
X$1695 145 146 147 251 148 252 257 258 cell_2rw
* cell instance $1696 r0 *1 23.5,92.69
X$1696 145 146 147 255 148 254 257 258 cell_2rw
* cell instance $1697 r0 *1 24.675,47.84
X$1697 149 150 151 199 152 201 257 258 cell_2rw
* cell instance $1698 m0 *1 24.675,50.83
X$1698 149 150 151 195 152 197 257 258 cell_2rw
* cell instance $1699 r0 *1 24.675,50.83
X$1699 149 150 151 202 152 194 257 258 cell_2rw
* cell instance $1700 m0 *1 24.675,53.82
X$1700 149 150 151 198 152 193 257 258 cell_2rw
* cell instance $1701 r0 *1 24.675,53.82
X$1701 149 150 151 196 152 200 257 258 cell_2rw
* cell instance $1702 m0 *1 24.675,56.81
X$1702 149 150 151 203 152 207 257 258 cell_2rw
* cell instance $1703 r0 *1 24.675,56.81
X$1703 149 150 151 206 152 208 257 258 cell_2rw
* cell instance $1704 m0 *1 24.675,59.8
X$1704 149 150 151 205 152 204 257 258 cell_2rw
* cell instance $1705 r0 *1 24.675,59.8
X$1705 149 150 151 214 152 213 257 258 cell_2rw
* cell instance $1706 m0 *1 24.675,62.79
X$1706 149 150 151 212 152 211 257 258 cell_2rw
* cell instance $1707 r0 *1 24.675,62.79
X$1707 149 150 151 210 152 209 257 258 cell_2rw
* cell instance $1708 m0 *1 24.675,65.78
X$1708 149 150 151 219 152 217 257 258 cell_2rw
* cell instance $1709 r0 *1 24.675,65.78
X$1709 149 150 151 216 152 215 257 258 cell_2rw
* cell instance $1710 m0 *1 24.675,68.77
X$1710 149 150 151 218 152 220 257 258 cell_2rw
* cell instance $1711 r0 *1 24.675,68.77
X$1711 149 150 151 224 152 223 257 258 cell_2rw
* cell instance $1712 m0 *1 24.675,71.76
X$1712 149 150 151 221 152 222 257 258 cell_2rw
* cell instance $1713 m0 *1 24.675,74.75
X$1713 149 150 151 231 152 232 257 258 cell_2rw
* cell instance $1714 r0 *1 24.675,71.76
X$1714 149 150 151 226 152 225 257 258 cell_2rw
* cell instance $1715 r0 *1 24.675,74.75
X$1715 149 150 151 230 152 229 257 258 cell_2rw
* cell instance $1716 m0 *1 24.675,77.74
X$1716 149 150 151 227 152 228 257 258 cell_2rw
* cell instance $1717 r0 *1 24.675,77.74
X$1717 149 150 151 237 152 238 257 258 cell_2rw
* cell instance $1718 m0 *1 24.675,80.73
X$1718 149 150 151 233 152 236 257 258 cell_2rw
* cell instance $1719 r0 *1 24.675,80.73
X$1719 149 150 151 235 152 234 257 258 cell_2rw
* cell instance $1720 m0 *1 24.675,83.72
X$1720 149 150 151 240 152 242 257 258 cell_2rw
* cell instance $1721 r0 *1 24.675,83.72
X$1721 149 150 151 239 152 241 257 258 cell_2rw
* cell instance $1722 m0 *1 24.675,86.71
X$1722 149 150 151 244 152 243 257 258 cell_2rw
* cell instance $1723 r0 *1 24.675,86.71
X$1723 149 150 151 245 152 247 257 258 cell_2rw
* cell instance $1724 m0 *1 24.675,89.7
X$1724 149 150 151 250 152 249 257 258 cell_2rw
* cell instance $1725 r0 *1 24.675,89.7
X$1725 149 150 151 246 152 248 257 258 cell_2rw
* cell instance $1726 m0 *1 24.675,92.69
X$1726 149 150 151 253 152 256 257 258 cell_2rw
* cell instance $1727 m0 *1 24.675,95.68
X$1727 149 150 151 251 152 252 257 258 cell_2rw
* cell instance $1728 r0 *1 24.675,92.69
X$1728 149 150 151 255 152 254 257 258 cell_2rw
* cell instance $1729 r0 *1 25.85,47.84
X$1729 153 154 155 199 156 201 257 258 cell_2rw
* cell instance $1730 m0 *1 25.85,50.83
X$1730 153 154 155 195 156 197 257 258 cell_2rw
* cell instance $1731 r0 *1 25.85,50.83
X$1731 153 154 155 202 156 194 257 258 cell_2rw
* cell instance $1732 m0 *1 25.85,53.82
X$1732 153 154 155 198 156 193 257 258 cell_2rw
* cell instance $1733 r0 *1 25.85,53.82
X$1733 153 154 155 196 156 200 257 258 cell_2rw
* cell instance $1734 m0 *1 25.85,56.81
X$1734 153 154 155 203 156 207 257 258 cell_2rw
* cell instance $1735 r0 *1 25.85,56.81
X$1735 153 154 155 206 156 208 257 258 cell_2rw
* cell instance $1736 m0 *1 25.85,59.8
X$1736 153 154 155 205 156 204 257 258 cell_2rw
* cell instance $1737 r0 *1 25.85,59.8
X$1737 153 154 155 214 156 213 257 258 cell_2rw
* cell instance $1738 m0 *1 25.85,62.79
X$1738 153 154 155 212 156 211 257 258 cell_2rw
* cell instance $1739 m0 *1 25.85,65.78
X$1739 153 154 155 219 156 217 257 258 cell_2rw
* cell instance $1740 r0 *1 25.85,62.79
X$1740 153 154 155 210 156 209 257 258 cell_2rw
* cell instance $1741 r0 *1 25.85,65.78
X$1741 153 154 155 216 156 215 257 258 cell_2rw
* cell instance $1742 m0 *1 25.85,68.77
X$1742 153 154 155 218 156 220 257 258 cell_2rw
* cell instance $1743 m0 *1 25.85,71.76
X$1743 153 154 155 221 156 222 257 258 cell_2rw
* cell instance $1744 r0 *1 25.85,68.77
X$1744 153 154 155 224 156 223 257 258 cell_2rw
* cell instance $1745 r0 *1 25.85,71.76
X$1745 153 154 155 226 156 225 257 258 cell_2rw
* cell instance $1746 m0 *1 25.85,74.75
X$1746 153 154 155 231 156 232 257 258 cell_2rw
* cell instance $1747 r0 *1 25.85,74.75
X$1747 153 154 155 230 156 229 257 258 cell_2rw
* cell instance $1748 m0 *1 25.85,77.74
X$1748 153 154 155 227 156 228 257 258 cell_2rw
* cell instance $1749 r0 *1 25.85,77.74
X$1749 153 154 155 237 156 238 257 258 cell_2rw
* cell instance $1750 m0 *1 25.85,80.73
X$1750 153 154 155 233 156 236 257 258 cell_2rw
* cell instance $1751 r0 *1 25.85,80.73
X$1751 153 154 155 235 156 234 257 258 cell_2rw
* cell instance $1752 m0 *1 25.85,83.72
X$1752 153 154 155 240 156 242 257 258 cell_2rw
* cell instance $1753 r0 *1 25.85,83.72
X$1753 153 154 155 239 156 241 257 258 cell_2rw
* cell instance $1754 m0 *1 25.85,86.71
X$1754 153 154 155 244 156 243 257 258 cell_2rw
* cell instance $1755 r0 *1 25.85,86.71
X$1755 153 154 155 245 156 247 257 258 cell_2rw
* cell instance $1756 m0 *1 25.85,89.7
X$1756 153 154 155 250 156 249 257 258 cell_2rw
* cell instance $1757 r0 *1 25.85,89.7
X$1757 153 154 155 246 156 248 257 258 cell_2rw
* cell instance $1758 m0 *1 25.85,92.69
X$1758 153 154 155 253 156 256 257 258 cell_2rw
* cell instance $1759 m0 *1 25.85,95.68
X$1759 153 154 155 251 156 252 257 258 cell_2rw
* cell instance $1760 r0 *1 25.85,92.69
X$1760 153 154 155 255 156 254 257 258 cell_2rw
* cell instance $1761 r0 *1 27.025,47.84
X$1761 157 158 159 199 160 201 257 258 cell_2rw
* cell instance $1762 m0 *1 27.025,50.83
X$1762 157 158 159 195 160 197 257 258 cell_2rw
* cell instance $1763 m0 *1 27.025,53.82
X$1763 157 158 159 198 160 193 257 258 cell_2rw
* cell instance $1764 r0 *1 27.025,50.83
X$1764 157 158 159 202 160 194 257 258 cell_2rw
* cell instance $1765 m0 *1 27.025,56.81
X$1765 157 158 159 203 160 207 257 258 cell_2rw
* cell instance $1766 r0 *1 27.025,53.82
X$1766 157 158 159 196 160 200 257 258 cell_2rw
* cell instance $1767 r0 *1 27.025,56.81
X$1767 157 158 159 206 160 208 257 258 cell_2rw
* cell instance $1768 m0 *1 27.025,59.8
X$1768 157 158 159 205 160 204 257 258 cell_2rw
* cell instance $1769 r0 *1 27.025,59.8
X$1769 157 158 159 214 160 213 257 258 cell_2rw
* cell instance $1770 m0 *1 27.025,62.79
X$1770 157 158 159 212 160 211 257 258 cell_2rw
* cell instance $1771 m0 *1 27.025,65.78
X$1771 157 158 159 219 160 217 257 258 cell_2rw
* cell instance $1772 r0 *1 27.025,62.79
X$1772 157 158 159 210 160 209 257 258 cell_2rw
* cell instance $1773 r0 *1 27.025,65.78
X$1773 157 158 159 216 160 215 257 258 cell_2rw
* cell instance $1774 m0 *1 27.025,68.77
X$1774 157 158 159 218 160 220 257 258 cell_2rw
* cell instance $1775 r0 *1 27.025,68.77
X$1775 157 158 159 224 160 223 257 258 cell_2rw
* cell instance $1776 m0 *1 27.025,71.76
X$1776 157 158 159 221 160 222 257 258 cell_2rw
* cell instance $1777 r0 *1 27.025,71.76
X$1777 157 158 159 226 160 225 257 258 cell_2rw
* cell instance $1778 m0 *1 27.025,74.75
X$1778 157 158 159 231 160 232 257 258 cell_2rw
* cell instance $1779 r0 *1 27.025,74.75
X$1779 157 158 159 230 160 229 257 258 cell_2rw
* cell instance $1780 m0 *1 27.025,77.74
X$1780 157 158 159 227 160 228 257 258 cell_2rw
* cell instance $1781 m0 *1 27.025,80.73
X$1781 157 158 159 233 160 236 257 258 cell_2rw
* cell instance $1782 r0 *1 27.025,77.74
X$1782 157 158 159 237 160 238 257 258 cell_2rw
* cell instance $1783 r0 *1 27.025,80.73
X$1783 157 158 159 235 160 234 257 258 cell_2rw
* cell instance $1784 m0 *1 27.025,83.72
X$1784 157 158 159 240 160 242 257 258 cell_2rw
* cell instance $1785 r0 *1 27.025,83.72
X$1785 157 158 159 239 160 241 257 258 cell_2rw
* cell instance $1786 m0 *1 27.025,86.71
X$1786 157 158 159 244 160 243 257 258 cell_2rw
* cell instance $1787 r0 *1 27.025,86.71
X$1787 157 158 159 245 160 247 257 258 cell_2rw
* cell instance $1788 m0 *1 27.025,89.7
X$1788 157 158 159 250 160 249 257 258 cell_2rw
* cell instance $1789 r0 *1 27.025,89.7
X$1789 157 158 159 246 160 248 257 258 cell_2rw
* cell instance $1790 m0 *1 27.025,92.69
X$1790 157 158 159 253 160 256 257 258 cell_2rw
* cell instance $1791 r0 *1 27.025,92.69
X$1791 157 158 159 255 160 254 257 258 cell_2rw
* cell instance $1792 m0 *1 27.025,95.68
X$1792 157 158 159 251 160 252 257 258 cell_2rw
* cell instance $1793 r0 *1 28.2,47.84
X$1793 161 162 163 199 164 201 257 258 cell_2rw
* cell instance $1794 m0 *1 28.2,50.83
X$1794 161 162 163 195 164 197 257 258 cell_2rw
* cell instance $1795 r0 *1 28.2,50.83
X$1795 161 162 163 202 164 194 257 258 cell_2rw
* cell instance $1796 m0 *1 28.2,53.82
X$1796 161 162 163 198 164 193 257 258 cell_2rw
* cell instance $1797 r0 *1 28.2,53.82
X$1797 161 162 163 196 164 200 257 258 cell_2rw
* cell instance $1798 m0 *1 28.2,56.81
X$1798 161 162 163 203 164 207 257 258 cell_2rw
* cell instance $1799 r0 *1 28.2,56.81
X$1799 161 162 163 206 164 208 257 258 cell_2rw
* cell instance $1800 m0 *1 28.2,59.8
X$1800 161 162 163 205 164 204 257 258 cell_2rw
* cell instance $1801 r0 *1 28.2,59.8
X$1801 161 162 163 214 164 213 257 258 cell_2rw
* cell instance $1802 m0 *1 28.2,62.79
X$1802 161 162 163 212 164 211 257 258 cell_2rw
* cell instance $1803 m0 *1 28.2,65.78
X$1803 161 162 163 219 164 217 257 258 cell_2rw
* cell instance $1804 r0 *1 28.2,62.79
X$1804 161 162 163 210 164 209 257 258 cell_2rw
* cell instance $1805 m0 *1 28.2,68.77
X$1805 161 162 163 218 164 220 257 258 cell_2rw
* cell instance $1806 r0 *1 28.2,65.78
X$1806 161 162 163 216 164 215 257 258 cell_2rw
* cell instance $1807 r0 *1 28.2,68.77
X$1807 161 162 163 224 164 223 257 258 cell_2rw
* cell instance $1808 m0 *1 28.2,71.76
X$1808 161 162 163 221 164 222 257 258 cell_2rw
* cell instance $1809 r0 *1 28.2,71.76
X$1809 161 162 163 226 164 225 257 258 cell_2rw
* cell instance $1810 m0 *1 28.2,74.75
X$1810 161 162 163 231 164 232 257 258 cell_2rw
* cell instance $1811 r0 *1 28.2,74.75
X$1811 161 162 163 230 164 229 257 258 cell_2rw
* cell instance $1812 m0 *1 28.2,77.74
X$1812 161 162 163 227 164 228 257 258 cell_2rw
* cell instance $1813 r0 *1 28.2,77.74
X$1813 161 162 163 237 164 238 257 258 cell_2rw
* cell instance $1814 m0 *1 28.2,80.73
X$1814 161 162 163 233 164 236 257 258 cell_2rw
* cell instance $1815 r0 *1 28.2,80.73
X$1815 161 162 163 235 164 234 257 258 cell_2rw
* cell instance $1816 m0 *1 28.2,83.72
X$1816 161 162 163 240 164 242 257 258 cell_2rw
* cell instance $1817 m0 *1 28.2,86.71
X$1817 161 162 163 244 164 243 257 258 cell_2rw
* cell instance $1818 r0 *1 28.2,83.72
X$1818 161 162 163 239 164 241 257 258 cell_2rw
* cell instance $1819 r0 *1 28.2,86.71
X$1819 161 162 163 245 164 247 257 258 cell_2rw
* cell instance $1820 m0 *1 28.2,89.7
X$1820 161 162 163 250 164 249 257 258 cell_2rw
* cell instance $1821 r0 *1 28.2,89.7
X$1821 161 162 163 246 164 248 257 258 cell_2rw
* cell instance $1822 m0 *1 28.2,92.69
X$1822 161 162 163 253 164 256 257 258 cell_2rw
* cell instance $1823 r0 *1 28.2,92.69
X$1823 161 162 163 255 164 254 257 258 cell_2rw
* cell instance $1824 m0 *1 28.2,95.68
X$1824 161 162 163 251 164 252 257 258 cell_2rw
* cell instance $1825 r0 *1 29.375,47.84
X$1825 165 166 167 199 168 201 257 258 cell_2rw
* cell instance $1826 m0 *1 29.375,50.83
X$1826 165 166 167 195 168 197 257 258 cell_2rw
* cell instance $1827 r0 *1 29.375,50.83
X$1827 165 166 167 202 168 194 257 258 cell_2rw
* cell instance $1828 m0 *1 29.375,53.82
X$1828 165 166 167 198 168 193 257 258 cell_2rw
* cell instance $1829 r0 *1 29.375,53.82
X$1829 165 166 167 196 168 200 257 258 cell_2rw
* cell instance $1830 m0 *1 29.375,56.81
X$1830 165 166 167 203 168 207 257 258 cell_2rw
* cell instance $1831 r0 *1 29.375,56.81
X$1831 165 166 167 206 168 208 257 258 cell_2rw
* cell instance $1832 m0 *1 29.375,59.8
X$1832 165 166 167 205 168 204 257 258 cell_2rw
* cell instance $1833 r0 *1 29.375,59.8
X$1833 165 166 167 214 168 213 257 258 cell_2rw
* cell instance $1834 m0 *1 29.375,62.79
X$1834 165 166 167 212 168 211 257 258 cell_2rw
* cell instance $1835 r0 *1 29.375,62.79
X$1835 165 166 167 210 168 209 257 258 cell_2rw
* cell instance $1836 m0 *1 29.375,65.78
X$1836 165 166 167 219 168 217 257 258 cell_2rw
* cell instance $1837 r0 *1 29.375,65.78
X$1837 165 166 167 216 168 215 257 258 cell_2rw
* cell instance $1838 m0 *1 29.375,68.77
X$1838 165 166 167 218 168 220 257 258 cell_2rw
* cell instance $1839 m0 *1 29.375,71.76
X$1839 165 166 167 221 168 222 257 258 cell_2rw
* cell instance $1840 r0 *1 29.375,68.77
X$1840 165 166 167 224 168 223 257 258 cell_2rw
* cell instance $1841 r0 *1 29.375,71.76
X$1841 165 166 167 226 168 225 257 258 cell_2rw
* cell instance $1842 m0 *1 29.375,74.75
X$1842 165 166 167 231 168 232 257 258 cell_2rw
* cell instance $1843 r0 *1 29.375,74.75
X$1843 165 166 167 230 168 229 257 258 cell_2rw
* cell instance $1844 m0 *1 29.375,77.74
X$1844 165 166 167 227 168 228 257 258 cell_2rw
* cell instance $1845 m0 *1 29.375,80.73
X$1845 165 166 167 233 168 236 257 258 cell_2rw
* cell instance $1846 r0 *1 29.375,77.74
X$1846 165 166 167 237 168 238 257 258 cell_2rw
* cell instance $1847 r0 *1 29.375,80.73
X$1847 165 166 167 235 168 234 257 258 cell_2rw
* cell instance $1848 m0 *1 29.375,83.72
X$1848 165 166 167 240 168 242 257 258 cell_2rw
* cell instance $1849 r0 *1 29.375,83.72
X$1849 165 166 167 239 168 241 257 258 cell_2rw
* cell instance $1850 m0 *1 29.375,86.71
X$1850 165 166 167 244 168 243 257 258 cell_2rw
* cell instance $1851 r0 *1 29.375,86.71
X$1851 165 166 167 245 168 247 257 258 cell_2rw
* cell instance $1852 m0 *1 29.375,89.7
X$1852 165 166 167 250 168 249 257 258 cell_2rw
* cell instance $1853 r0 *1 29.375,89.7
X$1853 165 166 167 246 168 248 257 258 cell_2rw
* cell instance $1854 m0 *1 29.375,92.69
X$1854 165 166 167 253 168 256 257 258 cell_2rw
* cell instance $1855 m0 *1 29.375,95.68
X$1855 165 166 167 251 168 252 257 258 cell_2rw
* cell instance $1856 r0 *1 29.375,92.69
X$1856 165 166 167 255 168 254 257 258 cell_2rw
* cell instance $1857 r0 *1 30.55,47.84
X$1857 169 170 171 199 172 201 257 258 cell_2rw
* cell instance $1858 m0 *1 30.55,50.83
X$1858 169 170 171 195 172 197 257 258 cell_2rw
* cell instance $1859 r0 *1 30.55,50.83
X$1859 169 170 171 202 172 194 257 258 cell_2rw
* cell instance $1860 m0 *1 30.55,53.82
X$1860 169 170 171 198 172 193 257 258 cell_2rw
* cell instance $1861 r0 *1 30.55,53.82
X$1861 169 170 171 196 172 200 257 258 cell_2rw
* cell instance $1862 m0 *1 30.55,56.81
X$1862 169 170 171 203 172 207 257 258 cell_2rw
* cell instance $1863 r0 *1 30.55,56.81
X$1863 169 170 171 206 172 208 257 258 cell_2rw
* cell instance $1864 m0 *1 30.55,59.8
X$1864 169 170 171 205 172 204 257 258 cell_2rw
* cell instance $1865 r0 *1 30.55,59.8
X$1865 169 170 171 214 172 213 257 258 cell_2rw
* cell instance $1866 m0 *1 30.55,62.79
X$1866 169 170 171 212 172 211 257 258 cell_2rw
* cell instance $1867 m0 *1 30.55,65.78
X$1867 169 170 171 219 172 217 257 258 cell_2rw
* cell instance $1868 r0 *1 30.55,62.79
X$1868 169 170 171 210 172 209 257 258 cell_2rw
* cell instance $1869 m0 *1 30.55,68.77
X$1869 169 170 171 218 172 220 257 258 cell_2rw
* cell instance $1870 r0 *1 30.55,65.78
X$1870 169 170 171 216 172 215 257 258 cell_2rw
* cell instance $1871 r0 *1 30.55,68.77
X$1871 169 170 171 224 172 223 257 258 cell_2rw
* cell instance $1872 m0 *1 30.55,71.76
X$1872 169 170 171 221 172 222 257 258 cell_2rw
* cell instance $1873 r0 *1 30.55,71.76
X$1873 169 170 171 226 172 225 257 258 cell_2rw
* cell instance $1874 m0 *1 30.55,74.75
X$1874 169 170 171 231 172 232 257 258 cell_2rw
* cell instance $1875 r0 *1 30.55,74.75
X$1875 169 170 171 230 172 229 257 258 cell_2rw
* cell instance $1876 m0 *1 30.55,77.74
X$1876 169 170 171 227 172 228 257 258 cell_2rw
* cell instance $1877 r0 *1 30.55,77.74
X$1877 169 170 171 237 172 238 257 258 cell_2rw
* cell instance $1878 m0 *1 30.55,80.73
X$1878 169 170 171 233 172 236 257 258 cell_2rw
* cell instance $1879 r0 *1 30.55,80.73
X$1879 169 170 171 235 172 234 257 258 cell_2rw
* cell instance $1880 m0 *1 30.55,83.72
X$1880 169 170 171 240 172 242 257 258 cell_2rw
* cell instance $1881 r0 *1 30.55,83.72
X$1881 169 170 171 239 172 241 257 258 cell_2rw
* cell instance $1882 m0 *1 30.55,86.71
X$1882 169 170 171 244 172 243 257 258 cell_2rw
* cell instance $1883 r0 *1 30.55,86.71
X$1883 169 170 171 245 172 247 257 258 cell_2rw
* cell instance $1884 m0 *1 30.55,89.7
X$1884 169 170 171 250 172 249 257 258 cell_2rw
* cell instance $1885 m0 *1 30.55,92.69
X$1885 169 170 171 253 172 256 257 258 cell_2rw
* cell instance $1886 r0 *1 30.55,89.7
X$1886 169 170 171 246 172 248 257 258 cell_2rw
* cell instance $1887 r0 *1 30.55,92.69
X$1887 169 170 171 255 172 254 257 258 cell_2rw
* cell instance $1888 m0 *1 30.55,95.68
X$1888 169 170 171 251 172 252 257 258 cell_2rw
* cell instance $1889 r0 *1 31.725,47.84
X$1889 173 174 175 199 176 201 257 258 cell_2rw
* cell instance $1890 m0 *1 31.725,50.83
X$1890 173 174 175 195 176 197 257 258 cell_2rw
* cell instance $1891 r0 *1 31.725,50.83
X$1891 173 174 175 202 176 194 257 258 cell_2rw
* cell instance $1892 m0 *1 31.725,53.82
X$1892 173 174 175 198 176 193 257 258 cell_2rw
* cell instance $1893 r0 *1 31.725,53.82
X$1893 173 174 175 196 176 200 257 258 cell_2rw
* cell instance $1894 m0 *1 31.725,56.81
X$1894 173 174 175 203 176 207 257 258 cell_2rw
* cell instance $1895 r0 *1 31.725,56.81
X$1895 173 174 175 206 176 208 257 258 cell_2rw
* cell instance $1896 m0 *1 31.725,59.8
X$1896 173 174 175 205 176 204 257 258 cell_2rw
* cell instance $1897 r0 *1 31.725,59.8
X$1897 173 174 175 214 176 213 257 258 cell_2rw
* cell instance $1898 m0 *1 31.725,62.79
X$1898 173 174 175 212 176 211 257 258 cell_2rw
* cell instance $1899 r0 *1 31.725,62.79
X$1899 173 174 175 210 176 209 257 258 cell_2rw
* cell instance $1900 m0 *1 31.725,65.78
X$1900 173 174 175 219 176 217 257 258 cell_2rw
* cell instance $1901 r0 *1 31.725,65.78
X$1901 173 174 175 216 176 215 257 258 cell_2rw
* cell instance $1902 m0 *1 31.725,68.77
X$1902 173 174 175 218 176 220 257 258 cell_2rw
* cell instance $1903 m0 *1 31.725,71.76
X$1903 173 174 175 221 176 222 257 258 cell_2rw
* cell instance $1904 r0 *1 31.725,68.77
X$1904 173 174 175 224 176 223 257 258 cell_2rw
* cell instance $1905 m0 *1 31.725,74.75
X$1905 173 174 175 231 176 232 257 258 cell_2rw
* cell instance $1906 r0 *1 31.725,71.76
X$1906 173 174 175 226 176 225 257 258 cell_2rw
* cell instance $1907 r0 *1 31.725,74.75
X$1907 173 174 175 230 176 229 257 258 cell_2rw
* cell instance $1908 m0 *1 31.725,77.74
X$1908 173 174 175 227 176 228 257 258 cell_2rw
* cell instance $1909 r0 *1 31.725,77.74
X$1909 173 174 175 237 176 238 257 258 cell_2rw
* cell instance $1910 m0 *1 31.725,80.73
X$1910 173 174 175 233 176 236 257 258 cell_2rw
* cell instance $1911 r0 *1 31.725,80.73
X$1911 173 174 175 235 176 234 257 258 cell_2rw
* cell instance $1912 m0 *1 31.725,83.72
X$1912 173 174 175 240 176 242 257 258 cell_2rw
* cell instance $1913 r0 *1 31.725,83.72
X$1913 173 174 175 239 176 241 257 258 cell_2rw
* cell instance $1914 m0 *1 31.725,86.71
X$1914 173 174 175 244 176 243 257 258 cell_2rw
* cell instance $1915 r0 *1 31.725,86.71
X$1915 173 174 175 245 176 247 257 258 cell_2rw
* cell instance $1916 m0 *1 31.725,89.7
X$1916 173 174 175 250 176 249 257 258 cell_2rw
* cell instance $1917 r0 *1 31.725,89.7
X$1917 173 174 175 246 176 248 257 258 cell_2rw
* cell instance $1918 m0 *1 31.725,92.69
X$1918 173 174 175 253 176 256 257 258 cell_2rw
* cell instance $1919 r0 *1 31.725,92.69
X$1919 173 174 175 255 176 254 257 258 cell_2rw
* cell instance $1920 m0 *1 31.725,95.68
X$1920 173 174 175 251 176 252 257 258 cell_2rw
* cell instance $1921 r0 *1 32.9,47.84
X$1921 177 178 179 199 180 201 257 258 cell_2rw
* cell instance $1922 m0 *1 32.9,50.83
X$1922 177 178 179 195 180 197 257 258 cell_2rw
* cell instance $1923 r0 *1 32.9,50.83
X$1923 177 178 179 202 180 194 257 258 cell_2rw
* cell instance $1924 m0 *1 32.9,53.82
X$1924 177 178 179 198 180 193 257 258 cell_2rw
* cell instance $1925 r0 *1 32.9,53.82
X$1925 177 178 179 196 180 200 257 258 cell_2rw
* cell instance $1926 m0 *1 32.9,56.81
X$1926 177 178 179 203 180 207 257 258 cell_2rw
* cell instance $1927 r0 *1 32.9,56.81
X$1927 177 178 179 206 180 208 257 258 cell_2rw
* cell instance $1928 m0 *1 32.9,59.8
X$1928 177 178 179 205 180 204 257 258 cell_2rw
* cell instance $1929 r0 *1 32.9,59.8
X$1929 177 178 179 214 180 213 257 258 cell_2rw
* cell instance $1930 m0 *1 32.9,62.79
X$1930 177 178 179 212 180 211 257 258 cell_2rw
* cell instance $1931 r0 *1 32.9,62.79
X$1931 177 178 179 210 180 209 257 258 cell_2rw
* cell instance $1932 m0 *1 32.9,65.78
X$1932 177 178 179 219 180 217 257 258 cell_2rw
* cell instance $1933 r0 *1 32.9,65.78
X$1933 177 178 179 216 180 215 257 258 cell_2rw
* cell instance $1934 m0 *1 32.9,68.77
X$1934 177 178 179 218 180 220 257 258 cell_2rw
* cell instance $1935 m0 *1 32.9,71.76
X$1935 177 178 179 221 180 222 257 258 cell_2rw
* cell instance $1936 r0 *1 32.9,68.77
X$1936 177 178 179 224 180 223 257 258 cell_2rw
* cell instance $1937 m0 *1 32.9,74.75
X$1937 177 178 179 231 180 232 257 258 cell_2rw
* cell instance $1938 r0 *1 32.9,71.76
X$1938 177 178 179 226 180 225 257 258 cell_2rw
* cell instance $1939 r0 *1 32.9,74.75
X$1939 177 178 179 230 180 229 257 258 cell_2rw
* cell instance $1940 m0 *1 32.9,77.74
X$1940 177 178 179 227 180 228 257 258 cell_2rw
* cell instance $1941 r0 *1 32.9,77.74
X$1941 177 178 179 237 180 238 257 258 cell_2rw
* cell instance $1942 m0 *1 32.9,80.73
X$1942 177 178 179 233 180 236 257 258 cell_2rw
* cell instance $1943 r0 *1 32.9,80.73
X$1943 177 178 179 235 180 234 257 258 cell_2rw
* cell instance $1944 m0 *1 32.9,83.72
X$1944 177 178 179 240 180 242 257 258 cell_2rw
* cell instance $1945 r0 *1 32.9,83.72
X$1945 177 178 179 239 180 241 257 258 cell_2rw
* cell instance $1946 m0 *1 32.9,86.71
X$1946 177 178 179 244 180 243 257 258 cell_2rw
* cell instance $1947 m0 *1 32.9,89.7
X$1947 177 178 179 250 180 249 257 258 cell_2rw
* cell instance $1948 r0 *1 32.9,86.71
X$1948 177 178 179 245 180 247 257 258 cell_2rw
* cell instance $1949 r0 *1 32.9,89.7
X$1949 177 178 179 246 180 248 257 258 cell_2rw
* cell instance $1950 m0 *1 32.9,92.69
X$1950 177 178 179 253 180 256 257 258 cell_2rw
* cell instance $1951 r0 *1 32.9,92.69
X$1951 177 178 179 255 180 254 257 258 cell_2rw
* cell instance $1952 m0 *1 32.9,95.68
X$1952 177 178 179 251 180 252 257 258 cell_2rw
* cell instance $1953 r0 *1 34.075,47.84
X$1953 181 182 183 199 184 201 257 258 cell_2rw
* cell instance $1954 m0 *1 34.075,50.83
X$1954 181 182 183 195 184 197 257 258 cell_2rw
* cell instance $1955 r0 *1 34.075,50.83
X$1955 181 182 183 202 184 194 257 258 cell_2rw
* cell instance $1956 m0 *1 34.075,53.82
X$1956 181 182 183 198 184 193 257 258 cell_2rw
* cell instance $1957 r0 *1 34.075,53.82
X$1957 181 182 183 196 184 200 257 258 cell_2rw
* cell instance $1958 m0 *1 34.075,56.81
X$1958 181 182 183 203 184 207 257 258 cell_2rw
* cell instance $1959 r0 *1 34.075,56.81
X$1959 181 182 183 206 184 208 257 258 cell_2rw
* cell instance $1960 m0 *1 34.075,59.8
X$1960 181 182 183 205 184 204 257 258 cell_2rw
* cell instance $1961 m0 *1 34.075,62.79
X$1961 181 182 183 212 184 211 257 258 cell_2rw
* cell instance $1962 r0 *1 34.075,59.8
X$1962 181 182 183 214 184 213 257 258 cell_2rw
* cell instance $1963 r0 *1 34.075,62.79
X$1963 181 182 183 210 184 209 257 258 cell_2rw
* cell instance $1964 m0 *1 34.075,65.78
X$1964 181 182 183 219 184 217 257 258 cell_2rw
* cell instance $1965 r0 *1 34.075,65.78
X$1965 181 182 183 216 184 215 257 258 cell_2rw
* cell instance $1966 m0 *1 34.075,68.77
X$1966 181 182 183 218 184 220 257 258 cell_2rw
* cell instance $1967 r0 *1 34.075,68.77
X$1967 181 182 183 224 184 223 257 258 cell_2rw
* cell instance $1968 m0 *1 34.075,71.76
X$1968 181 182 183 221 184 222 257 258 cell_2rw
* cell instance $1969 r0 *1 34.075,71.76
X$1969 181 182 183 226 184 225 257 258 cell_2rw
* cell instance $1970 m0 *1 34.075,74.75
X$1970 181 182 183 231 184 232 257 258 cell_2rw
* cell instance $1971 r0 *1 34.075,74.75
X$1971 181 182 183 230 184 229 257 258 cell_2rw
* cell instance $1972 m0 *1 34.075,77.74
X$1972 181 182 183 227 184 228 257 258 cell_2rw
* cell instance $1973 r0 *1 34.075,77.74
X$1973 181 182 183 237 184 238 257 258 cell_2rw
* cell instance $1974 m0 *1 34.075,80.73
X$1974 181 182 183 233 184 236 257 258 cell_2rw
* cell instance $1975 r0 *1 34.075,80.73
X$1975 181 182 183 235 184 234 257 258 cell_2rw
* cell instance $1976 m0 *1 34.075,83.72
X$1976 181 182 183 240 184 242 257 258 cell_2rw
* cell instance $1977 r0 *1 34.075,83.72
X$1977 181 182 183 239 184 241 257 258 cell_2rw
* cell instance $1978 m0 *1 34.075,86.71
X$1978 181 182 183 244 184 243 257 258 cell_2rw
* cell instance $1979 m0 *1 34.075,89.7
X$1979 181 182 183 250 184 249 257 258 cell_2rw
* cell instance $1980 r0 *1 34.075,86.71
X$1980 181 182 183 245 184 247 257 258 cell_2rw
* cell instance $1981 r0 *1 34.075,89.7
X$1981 181 182 183 246 184 248 257 258 cell_2rw
* cell instance $1982 m0 *1 34.075,92.69
X$1982 181 182 183 253 184 256 257 258 cell_2rw
* cell instance $1983 r0 *1 34.075,92.69
X$1983 181 182 183 255 184 254 257 258 cell_2rw
* cell instance $1984 m0 *1 34.075,95.68
X$1984 181 182 183 251 184 252 257 258 cell_2rw
* cell instance $1985 r0 *1 35.25,47.84
X$1985 185 186 187 199 188 201 257 258 cell_2rw
* cell instance $1986 m0 *1 35.25,50.83
X$1986 185 186 187 195 188 197 257 258 cell_2rw
* cell instance $1987 r0 *1 35.25,50.83
X$1987 185 186 187 202 188 194 257 258 cell_2rw
* cell instance $1988 m0 *1 35.25,53.82
X$1988 185 186 187 198 188 193 257 258 cell_2rw
* cell instance $1989 m0 *1 35.25,56.81
X$1989 185 186 187 203 188 207 257 258 cell_2rw
* cell instance $1990 r0 *1 35.25,53.82
X$1990 185 186 187 196 188 200 257 258 cell_2rw
* cell instance $1991 r0 *1 35.25,56.81
X$1991 185 186 187 206 188 208 257 258 cell_2rw
* cell instance $1992 m0 *1 35.25,59.8
X$1992 185 186 187 205 188 204 257 258 cell_2rw
* cell instance $1993 r0 *1 35.25,59.8
X$1993 185 186 187 214 188 213 257 258 cell_2rw
* cell instance $1994 m0 *1 35.25,62.79
X$1994 185 186 187 212 188 211 257 258 cell_2rw
* cell instance $1995 r0 *1 35.25,62.79
X$1995 185 186 187 210 188 209 257 258 cell_2rw
* cell instance $1996 m0 *1 35.25,65.78
X$1996 185 186 187 219 188 217 257 258 cell_2rw
* cell instance $1997 r0 *1 35.25,65.78
X$1997 185 186 187 216 188 215 257 258 cell_2rw
* cell instance $1998 m0 *1 35.25,68.77
X$1998 185 186 187 218 188 220 257 258 cell_2rw
* cell instance $1999 m0 *1 35.25,71.76
X$1999 185 186 187 221 188 222 257 258 cell_2rw
* cell instance $2000 r0 *1 35.25,68.77
X$2000 185 186 187 224 188 223 257 258 cell_2rw
* cell instance $2001 r0 *1 35.25,71.76
X$2001 185 186 187 226 188 225 257 258 cell_2rw
* cell instance $2002 m0 *1 35.25,74.75
X$2002 185 186 187 231 188 232 257 258 cell_2rw
* cell instance $2003 m0 *1 35.25,77.74
X$2003 185 186 187 227 188 228 257 258 cell_2rw
* cell instance $2004 r0 *1 35.25,74.75
X$2004 185 186 187 230 188 229 257 258 cell_2rw
* cell instance $2005 r0 *1 35.25,77.74
X$2005 185 186 187 237 188 238 257 258 cell_2rw
* cell instance $2006 m0 *1 35.25,80.73
X$2006 185 186 187 233 188 236 257 258 cell_2rw
* cell instance $2007 r0 *1 35.25,80.73
X$2007 185 186 187 235 188 234 257 258 cell_2rw
* cell instance $2008 m0 *1 35.25,83.72
X$2008 185 186 187 240 188 242 257 258 cell_2rw
* cell instance $2009 r0 *1 35.25,83.72
X$2009 185 186 187 239 188 241 257 258 cell_2rw
* cell instance $2010 m0 *1 35.25,86.71
X$2010 185 186 187 244 188 243 257 258 cell_2rw
* cell instance $2011 r0 *1 35.25,86.71
X$2011 185 186 187 245 188 247 257 258 cell_2rw
* cell instance $2012 m0 *1 35.25,89.7
X$2012 185 186 187 250 188 249 257 258 cell_2rw
* cell instance $2013 r0 *1 35.25,89.7
X$2013 185 186 187 246 188 248 257 258 cell_2rw
* cell instance $2014 m0 *1 35.25,92.69
X$2014 185 186 187 253 188 256 257 258 cell_2rw
* cell instance $2015 m0 *1 35.25,95.68
X$2015 185 186 187 251 188 252 257 258 cell_2rw
* cell instance $2016 r0 *1 35.25,92.69
X$2016 185 186 187 255 188 254 257 258 cell_2rw
* cell instance $2017 r0 *1 36.425,47.84
X$2017 189 190 191 199 192 201 257 258 cell_2rw
* cell instance $2018 m0 *1 36.425,50.83
X$2018 189 190 191 195 192 197 257 258 cell_2rw
* cell instance $2019 r0 *1 36.425,50.83
X$2019 189 190 191 202 192 194 257 258 cell_2rw
* cell instance $2020 m0 *1 36.425,53.82
X$2020 189 190 191 198 192 193 257 258 cell_2rw
* cell instance $2021 r0 *1 36.425,53.82
X$2021 189 190 191 196 192 200 257 258 cell_2rw
* cell instance $2022 m0 *1 36.425,56.81
X$2022 189 190 191 203 192 207 257 258 cell_2rw
* cell instance $2023 m0 *1 36.425,59.8
X$2023 189 190 191 205 192 204 257 258 cell_2rw
* cell instance $2024 r0 *1 36.425,56.81
X$2024 189 190 191 206 192 208 257 258 cell_2rw
* cell instance $2025 r0 *1 36.425,59.8
X$2025 189 190 191 214 192 213 257 258 cell_2rw
* cell instance $2026 m0 *1 36.425,62.79
X$2026 189 190 191 212 192 211 257 258 cell_2rw
* cell instance $2027 r0 *1 36.425,62.79
X$2027 189 190 191 210 192 209 257 258 cell_2rw
* cell instance $2028 m0 *1 36.425,65.78
X$2028 189 190 191 219 192 217 257 258 cell_2rw
* cell instance $2029 m0 *1 36.425,68.77
X$2029 189 190 191 218 192 220 257 258 cell_2rw
* cell instance $2030 r0 *1 36.425,65.78
X$2030 189 190 191 216 192 215 257 258 cell_2rw
* cell instance $2031 r0 *1 36.425,68.77
X$2031 189 190 191 224 192 223 257 258 cell_2rw
* cell instance $2032 m0 *1 36.425,71.76
X$2032 189 190 191 221 192 222 257 258 cell_2rw
* cell instance $2033 r0 *1 36.425,71.76
X$2033 189 190 191 226 192 225 257 258 cell_2rw
* cell instance $2034 m0 *1 36.425,74.75
X$2034 189 190 191 231 192 232 257 258 cell_2rw
* cell instance $2035 r0 *1 36.425,74.75
X$2035 189 190 191 230 192 229 257 258 cell_2rw
* cell instance $2036 m0 *1 36.425,77.74
X$2036 189 190 191 227 192 228 257 258 cell_2rw
* cell instance $2037 r0 *1 36.425,77.74
X$2037 189 190 191 237 192 238 257 258 cell_2rw
* cell instance $2038 m0 *1 36.425,80.73
X$2038 189 190 191 233 192 236 257 258 cell_2rw
* cell instance $2039 r0 *1 36.425,80.73
X$2039 189 190 191 235 192 234 257 258 cell_2rw
* cell instance $2040 m0 *1 36.425,83.72
X$2040 189 190 191 240 192 242 257 258 cell_2rw
* cell instance $2041 r0 *1 36.425,83.72
X$2041 189 190 191 239 192 241 257 258 cell_2rw
* cell instance $2042 m0 *1 36.425,86.71
X$2042 189 190 191 244 192 243 257 258 cell_2rw
* cell instance $2043 r0 *1 36.425,86.71
X$2043 189 190 191 245 192 247 257 258 cell_2rw
* cell instance $2044 m0 *1 36.425,89.7
X$2044 189 190 191 250 192 249 257 258 cell_2rw
* cell instance $2045 r0 *1 36.425,89.7
X$2045 189 190 191 246 192 248 257 258 cell_2rw
* cell instance $2046 m0 *1 36.425,92.69
X$2046 189 190 191 253 192 256 257 258 cell_2rw
* cell instance $2047 r0 *1 36.425,92.69
X$2047 189 190 191 255 192 254 257 258 cell_2rw
* cell instance $2048 m0 *1 36.425,95.68
X$2048 189 190 191 251 192 252 257 258 cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_bitcell_array_0

* cell custom_sram_1r1w_32_256_freepdk45_dummy_array
* pin wl_0_0
* pin wl_1_0
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_dummy_array 1 2 3 4
* net 1 wl_0_0
* net 2 wl_1_0
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 dummy_cell_2rw
* cell instance $2 r0 *1 1.175,0
X$2 2 1 3 4 dummy_cell_2rw
* cell instance $3 r0 *1 2.35,0
X$3 2 1 3 4 dummy_cell_2rw
* cell instance $4 r0 *1 3.525,0
X$4 2 1 3 4 dummy_cell_2rw
* cell instance $5 r0 *1 4.7,0
X$5 2 1 3 4 dummy_cell_2rw
* cell instance $6 r0 *1 5.875,0
X$6 2 1 3 4 dummy_cell_2rw
* cell instance $7 r0 *1 7.05,0
X$7 2 1 3 4 dummy_cell_2rw
* cell instance $8 r0 *1 8.225,0
X$8 2 1 3 4 dummy_cell_2rw
* cell instance $9 r0 *1 9.4,0
X$9 2 1 3 4 dummy_cell_2rw
* cell instance $10 r0 *1 10.575,0
X$10 2 1 3 4 dummy_cell_2rw
* cell instance $11 r0 *1 11.75,0
X$11 2 1 3 4 dummy_cell_2rw
* cell instance $12 r0 *1 12.925,0
X$12 2 1 3 4 dummy_cell_2rw
* cell instance $13 r0 *1 14.1,0
X$13 2 1 3 4 dummy_cell_2rw
* cell instance $14 r0 *1 15.275,0
X$14 2 1 3 4 dummy_cell_2rw
* cell instance $15 r0 *1 16.45,0
X$15 2 1 3 4 dummy_cell_2rw
* cell instance $16 r0 *1 17.625,0
X$16 2 1 3 4 dummy_cell_2rw
* cell instance $17 r0 *1 18.8,0
X$17 2 1 3 4 dummy_cell_2rw
* cell instance $18 r0 *1 19.975,0
X$18 2 1 3 4 dummy_cell_2rw
* cell instance $19 r0 *1 21.15,0
X$19 2 1 3 4 dummy_cell_2rw
* cell instance $20 r0 *1 22.325,0
X$20 2 1 3 4 dummy_cell_2rw
* cell instance $21 r0 *1 23.5,0
X$21 2 1 3 4 dummy_cell_2rw
* cell instance $22 r0 *1 24.675,0
X$22 2 1 3 4 dummy_cell_2rw
* cell instance $23 r0 *1 25.85,0
X$23 2 1 3 4 dummy_cell_2rw
* cell instance $24 r0 *1 27.025,0
X$24 2 1 3 4 dummy_cell_2rw
* cell instance $25 r0 *1 28.2,0
X$25 2 1 3 4 dummy_cell_2rw
* cell instance $26 r0 *1 29.375,0
X$26 2 1 3 4 dummy_cell_2rw
* cell instance $27 r0 *1 30.55,0
X$27 2 1 3 4 dummy_cell_2rw
* cell instance $28 r0 *1 31.725,0
X$28 2 1 3 4 dummy_cell_2rw
* cell instance $29 r0 *1 32.9,0
X$29 2 1 3 4 dummy_cell_2rw
* cell instance $30 r0 *1 34.075,0
X$30 2 1 3 4 dummy_cell_2rw
* cell instance $31 r0 *1 35.25,0
X$31 2 1 3 4 dummy_cell_2rw
* cell instance $32 r0 *1 36.425,0
X$32 2 1 3 4 dummy_cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_dummy_array

* cell custom_sram_1r1w_32_256_freepdk45_replica_column
* pin wl_0_0
* pin wl_1_0
* pin wl_1_1
* pin wl_0_1
* pin wl_0_2
* pin wl_1_2
* pin wl_1_3
* pin wl_0_3
* pin wl_0_4
* pin wl_1_4
* pin wl_1_5
* pin wl_0_5
* pin wl_0_6
* pin wl_1_6
* pin wl_1_7
* pin wl_0_7
* pin wl_0_8
* pin wl_1_8
* pin wl_1_9
* pin wl_0_9
* pin wl_0_10
* pin wl_1_10
* pin wl_1_11
* pin wl_0_11
* pin wl_0_12
* pin wl_1_12
* pin wl_1_13
* pin wl_0_13
* pin wl_0_14
* pin wl_1_14
* pin wl_1_15
* pin wl_0_15
* pin wl_0_16
* pin wl_1_16
* pin wl_1_17
* pin wl_0_17
* pin wl_0_18
* pin wl_1_18
* pin wl_1_19
* pin wl_0_19
* pin wl_0_20
* pin wl_1_20
* pin wl_1_21
* pin wl_0_21
* pin wl_0_22
* pin wl_1_22
* pin wl_1_23
* pin wl_0_23
* pin wl_0_24
* pin wl_1_24
* pin wl_1_25
* pin wl_0_25
* pin wl_0_26
* pin wl_1_26
* pin wl_1_27
* pin wl_0_27
* pin wl_0_28
* pin wl_1_28
* pin wl_1_29
* pin wl_0_29
* pin wl_0_30
* pin wl_1_30
* pin wl_1_31
* pin wl_0_31
* pin bl_0_0
* pin bl_1_0
* pin wl_0_32
* pin wl_1_32
* pin br_1_0
* pin br_0_0
* pin wl_1_33
* pin wl_0_33
* pin wl_0_34
* pin wl_1_34
* pin wl_1_35
* pin wl_0_35
* pin wl_0_36
* pin wl_1_36
* pin wl_1_37
* pin wl_0_37
* pin wl_0_38
* pin wl_1_38
* pin wl_1_39
* pin wl_0_39
* pin wl_0_40
* pin wl_1_40
* pin wl_1_41
* pin wl_0_41
* pin wl_0_42
* pin wl_1_42
* pin wl_1_43
* pin wl_0_43
* pin wl_0_44
* pin wl_1_44
* pin wl_1_45
* pin wl_0_45
* pin wl_0_46
* pin wl_1_46
* pin wl_1_47
* pin wl_0_47
* pin wl_0_48
* pin wl_1_48
* pin wl_1_49
* pin wl_0_49
* pin wl_0_50
* pin wl_1_50
* pin wl_1_51
* pin wl_0_51
* pin wl_0_52
* pin wl_1_52
* pin wl_1_53
* pin wl_0_53
* pin wl_0_54
* pin wl_1_54
* pin wl_1_55
* pin wl_0_55
* pin wl_0_56
* pin wl_1_56
* pin wl_1_57
* pin wl_0_57
* pin wl_0_58
* pin wl_1_58
* pin wl_1_59
* pin wl_0_59
* pin wl_0_60
* pin wl_1_60
* pin wl_1_61
* pin wl_0_61
* pin wl_0_62
* pin wl_1_62
* pin wl_1_63
* pin wl_0_63
* pin wl_0_64
* pin wl_1_64
* pin wl_1_65
* pin wl_0_65
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_replica_column 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36
+ 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129
+ 130 131 132 133 134 135 136 137 138
* net 1 wl_0_0
* net 2 wl_1_0
* net 3 wl_1_1
* net 4 wl_0_1
* net 5 wl_0_2
* net 6 wl_1_2
* net 7 wl_1_3
* net 8 wl_0_3
* net 9 wl_0_4
* net 10 wl_1_4
* net 11 wl_1_5
* net 12 wl_0_5
* net 13 wl_0_6
* net 14 wl_1_6
* net 15 wl_1_7
* net 16 wl_0_7
* net 17 wl_0_8
* net 18 wl_1_8
* net 19 wl_1_9
* net 20 wl_0_9
* net 21 wl_0_10
* net 22 wl_1_10
* net 23 wl_1_11
* net 24 wl_0_11
* net 25 wl_0_12
* net 26 wl_1_12
* net 27 wl_1_13
* net 28 wl_0_13
* net 29 wl_0_14
* net 30 wl_1_14
* net 31 wl_1_15
* net 32 wl_0_15
* net 33 wl_0_16
* net 34 wl_1_16
* net 35 wl_1_17
* net 36 wl_0_17
* net 37 wl_0_18
* net 38 wl_1_18
* net 39 wl_1_19
* net 40 wl_0_19
* net 41 wl_0_20
* net 42 wl_1_20
* net 43 wl_1_21
* net 44 wl_0_21
* net 45 wl_0_22
* net 46 wl_1_22
* net 47 wl_1_23
* net 48 wl_0_23
* net 49 wl_0_24
* net 50 wl_1_24
* net 51 wl_1_25
* net 52 wl_0_25
* net 53 wl_0_26
* net 54 wl_1_26
* net 55 wl_1_27
* net 56 wl_0_27
* net 57 wl_0_28
* net 58 wl_1_28
* net 59 wl_1_29
* net 60 wl_0_29
* net 61 wl_0_30
* net 62 wl_1_30
* net 63 wl_1_31
* net 64 wl_0_31
* net 65 bl_0_0
* net 66 bl_1_0
* net 67 wl_0_32
* net 68 wl_1_32
* net 69 br_1_0
* net 70 br_0_0
* net 71 wl_1_33
* net 72 wl_0_33
* net 73 wl_0_34
* net 74 wl_1_34
* net 75 wl_1_35
* net 76 wl_0_35
* net 77 wl_0_36
* net 78 wl_1_36
* net 79 wl_1_37
* net 80 wl_0_37
* net 81 wl_0_38
* net 82 wl_1_38
* net 83 wl_1_39
* net 84 wl_0_39
* net 85 wl_0_40
* net 86 wl_1_40
* net 87 wl_1_41
* net 88 wl_0_41
* net 89 wl_0_42
* net 90 wl_1_42
* net 91 wl_1_43
* net 92 wl_0_43
* net 93 wl_0_44
* net 94 wl_1_44
* net 95 wl_1_45
* net 96 wl_0_45
* net 97 wl_0_46
* net 98 wl_1_46
* net 99 wl_1_47
* net 100 wl_0_47
* net 101 wl_0_48
* net 102 wl_1_48
* net 103 wl_1_49
* net 104 wl_0_49
* net 105 wl_0_50
* net 106 wl_1_50
* net 107 wl_1_51
* net 108 wl_0_51
* net 109 wl_0_52
* net 110 wl_1_52
* net 111 wl_1_53
* net 112 wl_0_53
* net 113 wl_0_54
* net 114 wl_1_54
* net 115 wl_1_55
* net 116 wl_0_55
* net 117 wl_0_56
* net 118 wl_1_56
* net 119 wl_1_57
* net 120 wl_0_57
* net 121 wl_0_58
* net 122 wl_1_58
* net 123 wl_1_59
* net 124 wl_0_59
* net 125 wl_0_60
* net 126 wl_1_60
* net 127 wl_1_61
* net 128 wl_0_61
* net 129 wl_0_62
* net 130 wl_1_62
* net 131 wl_1_63
* net 132 wl_0_63
* net 133 wl_0_64
* net 134 wl_1_64
* net 135 wl_1_65
* net 136 wl_0_65
* net 137 vdd
* net 138 gnd
* cell instance $1 m0 *1 0,1.495
X$1 65 66 69 2 70 1 137 138 replica_cell_2rw
* cell instance $2 r0 *1 0,1.495
X$2 65 66 69 3 70 4 137 138 replica_cell_2rw
* cell instance $3 m0 *1 0,4.485
X$3 65 66 69 6 70 5 137 138 replica_cell_2rw
* cell instance $4 r0 *1 0,4.485
X$4 65 66 69 7 70 8 137 138 replica_cell_2rw
* cell instance $5 m0 *1 0,7.475
X$5 65 66 69 10 70 9 137 138 replica_cell_2rw
* cell instance $6 r0 *1 0,7.475
X$6 65 66 69 11 70 12 137 138 replica_cell_2rw
* cell instance $7 m0 *1 0,10.465
X$7 65 66 69 14 70 13 137 138 replica_cell_2rw
* cell instance $8 r0 *1 0,10.465
X$8 65 66 69 15 70 16 137 138 replica_cell_2rw
* cell instance $9 m0 *1 0,13.455
X$9 65 66 69 18 70 17 137 138 replica_cell_2rw
* cell instance $10 r0 *1 0,13.455
X$10 65 66 69 19 70 20 137 138 replica_cell_2rw
* cell instance $11 m0 *1 0,16.445
X$11 65 66 69 22 70 21 137 138 replica_cell_2rw
* cell instance $12 r0 *1 0,16.445
X$12 65 66 69 23 70 24 137 138 replica_cell_2rw
* cell instance $13 m0 *1 0,19.435
X$13 65 66 69 26 70 25 137 138 replica_cell_2rw
* cell instance $14 r0 *1 0,19.435
X$14 65 66 69 27 70 28 137 138 replica_cell_2rw
* cell instance $15 m0 *1 0,22.425
X$15 65 66 69 30 70 29 137 138 replica_cell_2rw
* cell instance $16 r0 *1 0,22.425
X$16 65 66 69 31 70 32 137 138 replica_cell_2rw
* cell instance $17 m0 *1 0,25.415
X$17 65 66 69 34 70 33 137 138 replica_cell_2rw
* cell instance $18 r0 *1 0,25.415
X$18 65 66 69 35 70 36 137 138 replica_cell_2rw
* cell instance $19 m0 *1 0,28.405
X$19 65 66 69 38 70 37 137 138 replica_cell_2rw
* cell instance $20 r0 *1 0,28.405
X$20 65 66 69 39 70 40 137 138 replica_cell_2rw
* cell instance $21 m0 *1 0,31.395
X$21 65 66 69 42 70 41 137 138 replica_cell_2rw
* cell instance $22 r0 *1 0,31.395
X$22 65 66 69 43 70 44 137 138 replica_cell_2rw
* cell instance $23 m0 *1 0,34.385
X$23 65 66 69 46 70 45 137 138 replica_cell_2rw
* cell instance $24 r0 *1 0,34.385
X$24 65 66 69 47 70 48 137 138 replica_cell_2rw
* cell instance $25 m0 *1 0,37.375
X$25 65 66 69 50 70 49 137 138 replica_cell_2rw
* cell instance $26 r0 *1 0,37.375
X$26 65 66 69 51 70 52 137 138 replica_cell_2rw
* cell instance $27 m0 *1 0,40.365
X$27 65 66 69 54 70 53 137 138 replica_cell_2rw
* cell instance $28 r0 *1 0,40.365
X$28 65 66 69 55 70 56 137 138 replica_cell_2rw
* cell instance $29 m0 *1 0,43.355
X$29 65 66 69 58 70 57 137 138 replica_cell_2rw
* cell instance $30 r0 *1 0,43.355
X$30 65 66 69 59 70 60 137 138 replica_cell_2rw
* cell instance $31 m0 *1 0,46.345
X$31 65 66 69 62 70 61 137 138 replica_cell_2rw
* cell instance $32 r0 *1 0,46.345
X$32 65 66 69 63 70 64 137 138 replica_cell_2rw
* cell instance $33 m0 *1 0,49.335
X$33 65 66 69 68 70 67 137 138 replica_cell_2rw
* cell instance $34 r0 *1 0,49.335
X$34 65 66 69 71 70 72 137 138 replica_cell_2rw
* cell instance $35 m0 *1 0,52.325
X$35 65 66 69 74 70 73 137 138 replica_cell_2rw
* cell instance $36 r0 *1 0,52.325
X$36 65 66 69 75 70 76 137 138 replica_cell_2rw
* cell instance $37 m0 *1 0,55.315
X$37 65 66 69 78 70 77 137 138 replica_cell_2rw
* cell instance $38 r0 *1 0,55.315
X$38 65 66 69 79 70 80 137 138 replica_cell_2rw
* cell instance $39 m0 *1 0,58.305
X$39 65 66 69 82 70 81 137 138 replica_cell_2rw
* cell instance $40 r0 *1 0,58.305
X$40 65 66 69 83 70 84 137 138 replica_cell_2rw
* cell instance $41 m0 *1 0,61.295
X$41 65 66 69 86 70 85 137 138 replica_cell_2rw
* cell instance $42 r0 *1 0,61.295
X$42 65 66 69 87 70 88 137 138 replica_cell_2rw
* cell instance $43 m0 *1 0,64.285
X$43 65 66 69 90 70 89 137 138 replica_cell_2rw
* cell instance $44 r0 *1 0,64.285
X$44 65 66 69 91 70 92 137 138 replica_cell_2rw
* cell instance $45 m0 *1 0,67.275
X$45 65 66 69 94 70 93 137 138 replica_cell_2rw
* cell instance $46 r0 *1 0,67.275
X$46 65 66 69 95 70 96 137 138 replica_cell_2rw
* cell instance $47 m0 *1 0,70.265
X$47 65 66 69 98 70 97 137 138 replica_cell_2rw
* cell instance $48 r0 *1 0,70.265
X$48 65 66 69 99 70 100 137 138 replica_cell_2rw
* cell instance $49 m0 *1 0,73.255
X$49 65 66 69 102 70 101 137 138 replica_cell_2rw
* cell instance $50 r0 *1 0,73.255
X$50 65 66 69 103 70 104 137 138 replica_cell_2rw
* cell instance $51 m0 *1 0,76.245
X$51 65 66 69 106 70 105 137 138 replica_cell_2rw
* cell instance $52 r0 *1 0,76.245
X$52 65 66 69 107 70 108 137 138 replica_cell_2rw
* cell instance $53 m0 *1 0,79.235
X$53 65 66 69 110 70 109 137 138 replica_cell_2rw
* cell instance $54 r0 *1 0,79.235
X$54 65 66 69 111 70 112 137 138 replica_cell_2rw
* cell instance $55 m0 *1 0,82.225
X$55 65 66 69 114 70 113 137 138 replica_cell_2rw
* cell instance $56 r0 *1 0,82.225
X$56 65 66 69 115 70 116 137 138 replica_cell_2rw
* cell instance $57 m0 *1 0,85.215
X$57 65 66 69 118 70 117 137 138 replica_cell_2rw
* cell instance $58 r0 *1 0,85.215
X$58 65 66 69 119 70 120 137 138 replica_cell_2rw
* cell instance $59 m0 *1 0,88.205
X$59 65 66 69 122 70 121 137 138 replica_cell_2rw
* cell instance $60 r0 *1 0,88.205
X$60 65 66 69 123 70 124 137 138 replica_cell_2rw
* cell instance $61 m0 *1 0,91.195
X$61 65 66 69 126 70 125 137 138 replica_cell_2rw
* cell instance $62 r0 *1 0,91.195
X$62 65 66 69 127 70 128 137 138 replica_cell_2rw
* cell instance $63 m0 *1 0,94.185
X$63 65 66 69 130 70 129 137 138 replica_cell_2rw
* cell instance $64 r0 *1 0,94.185
X$64 65 66 69 131 70 132 137 138 replica_cell_2rw
* cell instance $65 m0 *1 0,97.175
X$65 65 66 69 134 70 133 137 138 replica_cell_2rw
* cell instance $66 r0 *1 0,97.175
X$66 135 136 137 138 dummy_cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_replica_column

* cell custom_sram_1r1w_32_256_freepdk45_bitcell_array
* pin wl_0_2
* pin wl_1_2
* pin wl_0_1
* pin wl_1_1
* pin wl_0_0
* pin wl_1_0
* pin wl_1_4
* pin wl_0_5
* pin wl_1_5
* pin wl_0_4
* pin wl_1_3
* pin wl_0_3
* pin wl_1_7
* pin wl_0_7
* pin wl_0_8
* pin wl_1_8
* pin wl_1_6
* pin wl_0_6
* pin wl_0_10
* pin wl_1_10
* pin wl_1_11
* pin wl_0_11
* pin wl_0_9
* pin wl_1_9
* pin wl_0_14
* pin wl_1_13
* pin wl_1_12
* pin wl_1_14
* pin wl_0_13
* pin wl_0_12
* pin wl_1_16
* pin wl_0_17
* pin wl_0_16
* pin wl_1_17
* pin wl_1_15
* pin wl_0_15
* pin wl_1_20
* pin wl_0_20
* pin wl_0_18
* pin wl_0_19
* pin wl_1_19
* pin wl_1_18
* pin wl_0_22
* pin wl_1_22
* pin wl_1_23
* pin wl_0_23
* pin wl_0_21
* pin wl_1_21
* pin wl_0_25
* pin wl_0_26
* pin wl_1_26
* pin wl_0_24
* pin wl_1_24
* pin wl_1_25
* pin wl_0_28
* pin wl_1_28
* pin wl_0_29
* pin wl_0_27
* pin wl_1_27
* pin wl_1_29
* pin bl_0_0
* pin bl_1_0
* pin br_1_0
* pin br_0_0
* pin bl_0_1
* pin bl_1_1
* pin br_1_1
* pin br_0_1
* pin bl_0_2
* pin bl_1_2
* pin br_1_2
* pin br_0_2
* pin bl_0_3
* pin bl_1_3
* pin br_1_3
* pin br_0_3
* pin bl_0_4
* pin bl_1_4
* pin br_1_4
* pin br_0_4
* pin bl_0_5
* pin bl_1_5
* pin br_1_5
* pin br_0_5
* pin bl_0_6
* pin bl_1_6
* pin br_1_6
* pin br_0_6
* pin bl_0_7
* pin bl_1_7
* pin br_1_7
* pin br_0_7
* pin bl_0_8
* pin bl_1_8
* pin br_1_8
* pin br_0_8
* pin bl_0_9
* pin bl_1_9
* pin br_1_9
* pin br_0_9
* pin bl_0_10
* pin bl_1_10
* pin br_1_10
* pin br_0_10
* pin bl_0_11
* pin bl_1_11
* pin br_1_11
* pin br_0_11
* pin bl_0_12
* pin bl_1_12
* pin br_1_12
* pin br_0_12
* pin bl_0_13
* pin bl_1_13
* pin br_1_13
* pin br_0_13
* pin bl_0_14
* pin bl_1_14
* pin br_1_14
* pin br_0_14
* pin bl_0_15
* pin bl_1_15
* pin br_1_15
* pin br_0_15
* pin wl_0_31
* pin wl_1_31
* pin wl_1_30
* pin wl_0_30
* pin bl_0_16
* pin bl_1_16
* pin br_1_16
* pin br_0_16
* pin bl_0_17
* pin bl_1_17
* pin br_1_17
* pin br_0_17
* pin bl_0_18
* pin bl_1_18
* pin br_1_18
* pin br_0_18
* pin bl_0_19
* pin bl_1_19
* pin br_1_19
* pin br_0_19
* pin bl_0_20
* pin bl_1_20
* pin br_1_20
* pin br_0_20
* pin bl_0_21
* pin bl_1_21
* pin br_1_21
* pin br_0_21
* pin bl_0_22
* pin bl_1_22
* pin br_1_22
* pin br_0_22
* pin bl_0_23
* pin bl_1_23
* pin br_1_23
* pin br_0_23
* pin bl_0_24
* pin bl_1_24
* pin br_1_24
* pin br_0_24
* pin bl_0_25
* pin bl_1_25
* pin br_1_25
* pin br_0_25
* pin bl_0_26
* pin bl_1_26
* pin br_1_26
* pin br_0_26
* pin bl_0_27
* pin bl_1_27
* pin br_1_27
* pin br_0_27
* pin bl_0_28
* pin bl_1_28
* pin br_1_28
* pin br_0_28
* pin bl_0_29
* pin bl_1_29
* pin br_1_29
* pin br_0_29
* pin bl_0_30
* pin bl_1_30
* pin br_1_30
* pin br_0_30
* pin bl_0_31
* pin bl_1_31
* pin br_1_31
* pin br_0_31
* pin wl_0_35
* pin wl_0_34
* pin wl_1_33
* pin wl_1_36
* pin wl_0_33
* pin wl_1_35
* pin wl_1_32
* pin wl_0_36
* pin wl_0_32
* pin wl_1_34
* pin wl_1_37
* pin wl_0_39
* pin wl_1_39
* pin wl_1_38
* pin wl_0_37
* pin wl_0_38
* pin wl_0_42
* pin wl_1_42
* pin wl_0_41
* pin wl_1_41
* pin wl_0_40
* pin wl_1_40
* pin wl_0_44
* pin wl_1_44
* pin wl_0_43
* pin wl_1_45
* pin wl_1_43
* pin wl_0_45
* pin wl_1_47
* pin wl_0_47
* pin wl_0_46
* pin wl_1_46
* pin wl_0_48
* pin wl_1_48
* pin wl_1_51
* pin wl_0_51
* pin wl_0_50
* pin wl_1_50
* pin wl_1_49
* pin wl_0_49
* pin wl_1_53
* pin wl_0_54
* pin wl_1_54
* pin wl_0_53
* pin wl_1_52
* pin wl_0_52
* pin wl_1_56
* pin wl_1_55
* pin wl_0_56
* pin wl_0_55
* pin wl_0_57
* pin wl_1_57
* pin wl_1_58
* pin wl_1_60
* pin wl_0_58
* pin wl_0_60
* pin wl_0_59
* pin wl_1_59
* pin wl_1_63
* pin wl_0_63
* pin wl_1_61
* pin wl_0_62
* pin wl_1_62
* pin wl_0_61
* pin vdd
* pin gnd
.SUBCKT custom_sram_1r1w_32_256_freepdk45_bitcell_array 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37
+ 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89
+ 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111
+ 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130
+ 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149
+ 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168
+ 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187
+ 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206
+ 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225
+ 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244
+ 245 246 247 248 249 250 251 252 253 254 255 256 257 258
* net 1 wl_0_2
* net 2 wl_1_2
* net 3 wl_0_1
* net 4 wl_1_1
* net 5 wl_0_0
* net 6 wl_1_0
* net 7 wl_1_4
* net 8 wl_0_5
* net 9 wl_1_5
* net 10 wl_0_4
* net 11 wl_1_3
* net 12 wl_0_3
* net 13 wl_1_7
* net 14 wl_0_7
* net 15 wl_0_8
* net 16 wl_1_8
* net 17 wl_1_6
* net 18 wl_0_6
* net 19 wl_0_10
* net 20 wl_1_10
* net 21 wl_1_11
* net 22 wl_0_11
* net 23 wl_0_9
* net 24 wl_1_9
* net 25 wl_0_14
* net 26 wl_1_13
* net 27 wl_1_12
* net 28 wl_1_14
* net 29 wl_0_13
* net 30 wl_0_12
* net 31 wl_1_16
* net 32 wl_0_17
* net 33 wl_0_16
* net 34 wl_1_17
* net 35 wl_1_15
* net 36 wl_0_15
* net 37 wl_1_20
* net 38 wl_0_20
* net 39 wl_0_18
* net 40 wl_0_19
* net 41 wl_1_19
* net 42 wl_1_18
* net 43 wl_0_22
* net 44 wl_1_22
* net 45 wl_1_23
* net 46 wl_0_23
* net 47 wl_0_21
* net 48 wl_1_21
* net 49 wl_0_25
* net 50 wl_0_26
* net 51 wl_1_26
* net 52 wl_0_24
* net 53 wl_1_24
* net 54 wl_1_25
* net 55 wl_0_28
* net 56 wl_1_28
* net 57 wl_0_29
* net 58 wl_0_27
* net 59 wl_1_27
* net 60 wl_1_29
* net 61 bl_0_0
* net 62 bl_1_0
* net 63 br_1_0
* net 64 br_0_0
* net 65 bl_0_1
* net 66 bl_1_1
* net 67 br_1_1
* net 68 br_0_1
* net 69 bl_0_2
* net 70 bl_1_2
* net 71 br_1_2
* net 72 br_0_2
* net 73 bl_0_3
* net 74 bl_1_3
* net 75 br_1_3
* net 76 br_0_3
* net 77 bl_0_4
* net 78 bl_1_4
* net 79 br_1_4
* net 80 br_0_4
* net 81 bl_0_5
* net 82 bl_1_5
* net 83 br_1_5
* net 84 br_0_5
* net 85 bl_0_6
* net 86 bl_1_6
* net 87 br_1_6
* net 88 br_0_6
* net 89 bl_0_7
* net 90 bl_1_7
* net 91 br_1_7
* net 92 br_0_7
* net 93 bl_0_8
* net 94 bl_1_8
* net 95 br_1_8
* net 96 br_0_8
* net 97 bl_0_9
* net 98 bl_1_9
* net 99 br_1_9
* net 100 br_0_9
* net 101 bl_0_10
* net 102 bl_1_10
* net 103 br_1_10
* net 104 br_0_10
* net 105 bl_0_11
* net 106 bl_1_11
* net 107 br_1_11
* net 108 br_0_11
* net 109 bl_0_12
* net 110 bl_1_12
* net 111 br_1_12
* net 112 br_0_12
* net 113 bl_0_13
* net 114 bl_1_13
* net 115 br_1_13
* net 116 br_0_13
* net 117 bl_0_14
* net 118 bl_1_14
* net 119 br_1_14
* net 120 br_0_14
* net 121 bl_0_15
* net 122 bl_1_15
* net 123 br_1_15
* net 124 br_0_15
* net 125 wl_0_31
* net 126 wl_1_31
* net 127 wl_1_30
* net 128 wl_0_30
* net 129 bl_0_16
* net 130 bl_1_16
* net 131 br_1_16
* net 132 br_0_16
* net 133 bl_0_17
* net 134 bl_1_17
* net 135 br_1_17
* net 136 br_0_17
* net 137 bl_0_18
* net 138 bl_1_18
* net 139 br_1_18
* net 140 br_0_18
* net 141 bl_0_19
* net 142 bl_1_19
* net 143 br_1_19
* net 144 br_0_19
* net 145 bl_0_20
* net 146 bl_1_20
* net 147 br_1_20
* net 148 br_0_20
* net 149 bl_0_21
* net 150 bl_1_21
* net 151 br_1_21
* net 152 br_0_21
* net 153 bl_0_22
* net 154 bl_1_22
* net 155 br_1_22
* net 156 br_0_22
* net 157 bl_0_23
* net 158 bl_1_23
* net 159 br_1_23
* net 160 br_0_23
* net 161 bl_0_24
* net 162 bl_1_24
* net 163 br_1_24
* net 164 br_0_24
* net 165 bl_0_25
* net 166 bl_1_25
* net 167 br_1_25
* net 168 br_0_25
* net 169 bl_0_26
* net 170 bl_1_26
* net 171 br_1_26
* net 172 br_0_26
* net 173 bl_0_27
* net 174 bl_1_27
* net 175 br_1_27
* net 176 br_0_27
* net 177 bl_0_28
* net 178 bl_1_28
* net 179 br_1_28
* net 180 br_0_28
* net 181 bl_0_29
* net 182 bl_1_29
* net 183 br_1_29
* net 184 br_0_29
* net 185 bl_0_30
* net 186 bl_1_30
* net 187 br_1_30
* net 188 br_0_30
* net 189 bl_0_31
* net 190 bl_1_31
* net 191 br_1_31
* net 192 br_0_31
* net 193 wl_0_35
* net 194 wl_0_34
* net 195 wl_1_33
* net 196 wl_1_36
* net 197 wl_0_33
* net 198 wl_1_35
* net 199 wl_1_32
* net 200 wl_0_36
* net 201 wl_0_32
* net 202 wl_1_34
* net 203 wl_1_37
* net 204 wl_0_39
* net 205 wl_1_39
* net 206 wl_1_38
* net 207 wl_0_37
* net 208 wl_0_38
* net 209 wl_0_42
* net 210 wl_1_42
* net 211 wl_0_41
* net 212 wl_1_41
* net 213 wl_0_40
* net 214 wl_1_40
* net 215 wl_0_44
* net 216 wl_1_44
* net 217 wl_0_43
* net 218 wl_1_45
* net 219 wl_1_43
* net 220 wl_0_45
* net 221 wl_1_47
* net 222 wl_0_47
* net 223 wl_0_46
* net 224 wl_1_46
* net 225 wl_0_48
* net 226 wl_1_48
* net 227 wl_1_51
* net 228 wl_0_51
* net 229 wl_0_50
* net 230 wl_1_50
* net 231 wl_1_49
* net 232 wl_0_49
* net 233 wl_1_53
* net 234 wl_0_54
* net 235 wl_1_54
* net 236 wl_0_53
* net 237 wl_1_52
* net 238 wl_0_52
* net 239 wl_1_56
* net 240 wl_1_55
* net 241 wl_0_56
* net 242 wl_0_55
* net 243 wl_0_57
* net 244 wl_1_57
* net 245 wl_1_58
* net 246 wl_1_60
* net 247 wl_0_58
* net 248 wl_0_60
* net 249 wl_0_59
* net 250 wl_1_59
* net 251 wl_1_63
* net 252 wl_0_63
* net 253 wl_1_61
* net 254 wl_0_62
* net 255 wl_1_62
* net 256 wl_0_61
* net 257 vdd
* net 258 gnd
* cell instance $1 r0 *1 1.175,2.99
X$1 65 66 67 2 68 1 257 258 cell_2rw
* cell instance $2 r0 *1 0,2.99
X$2 61 62 63 2 64 1 257 258 cell_2rw
* cell instance $3 r0 *1 2.35,2.99
X$3 69 70 71 2 72 1 257 258 cell_2rw
* cell instance $4 r0 *1 3.525,2.99
X$4 73 74 75 2 76 1 257 258 cell_2rw
* cell instance $5 r0 *1 4.7,2.99
X$5 77 78 79 2 80 1 257 258 cell_2rw
* cell instance $6 r0 *1 5.875,2.99
X$6 81 82 83 2 84 1 257 258 cell_2rw
* cell instance $7 r0 *1 7.05,2.99
X$7 85 86 87 2 88 1 257 258 cell_2rw
* cell instance $8 r0 *1 8.225,2.99
X$8 89 90 91 2 92 1 257 258 cell_2rw
* cell instance $9 r0 *1 9.4,2.99
X$9 93 94 95 2 96 1 257 258 cell_2rw
* cell instance $10 r0 *1 10.575,2.99
X$10 97 98 99 2 100 1 257 258 cell_2rw
* cell instance $11 r0 *1 11.75,2.99
X$11 101 102 103 2 104 1 257 258 cell_2rw
* cell instance $12 r0 *1 12.925,2.99
X$12 105 106 107 2 108 1 257 258 cell_2rw
* cell instance $13 r0 *1 14.1,2.99
X$13 109 110 111 2 112 1 257 258 cell_2rw
* cell instance $14 r0 *1 15.275,2.99
X$14 113 114 115 2 116 1 257 258 cell_2rw
* cell instance $15 r0 *1 16.45,2.99
X$15 117 118 119 2 120 1 257 258 cell_2rw
* cell instance $16 r0 *1 17.625,2.99
X$16 121 122 123 2 124 1 257 258 cell_2rw
* cell instance $17 r0 *1 18.8,2.99
X$17 129 130 131 2 132 1 257 258 cell_2rw
* cell instance $18 r0 *1 19.975,2.99
X$18 133 134 135 2 136 1 257 258 cell_2rw
* cell instance $19 r0 *1 21.15,2.99
X$19 137 138 139 2 140 1 257 258 cell_2rw
* cell instance $20 r0 *1 22.325,2.99
X$20 141 142 143 2 144 1 257 258 cell_2rw
* cell instance $21 r0 *1 23.5,2.99
X$21 145 146 147 2 148 1 257 258 cell_2rw
* cell instance $22 r0 *1 24.675,2.99
X$22 149 150 151 2 152 1 257 258 cell_2rw
* cell instance $23 r0 *1 25.85,2.99
X$23 153 154 155 2 156 1 257 258 cell_2rw
* cell instance $24 r0 *1 27.025,2.99
X$24 157 158 159 2 160 1 257 258 cell_2rw
* cell instance $25 r0 *1 28.2,2.99
X$25 161 162 163 2 164 1 257 258 cell_2rw
* cell instance $26 r0 *1 29.375,2.99
X$26 165 166 167 2 168 1 257 258 cell_2rw
* cell instance $27 r0 *1 30.55,2.99
X$27 169 170 171 2 172 1 257 258 cell_2rw
* cell instance $28 r0 *1 31.725,2.99
X$28 173 174 175 2 176 1 257 258 cell_2rw
* cell instance $29 r0 *1 32.9,2.99
X$29 177 178 179 2 180 1 257 258 cell_2rw
* cell instance $30 r0 *1 34.075,2.99
X$30 181 182 183 2 184 1 257 258 cell_2rw
* cell instance $31 r0 *1 35.25,2.99
X$31 185 186 187 2 188 1 257 258 cell_2rw
* cell instance $32 r0 *1 36.425,2.99
X$32 189 190 191 2 192 1 257 258 cell_2rw
* cell instance $33 m0 *1 1.175,2.99
X$33 65 66 67 4 68 3 257 258 cell_2rw
* cell instance $34 m0 *1 0,2.99
X$34 61 62 63 4 64 3 257 258 cell_2rw
* cell instance $35 m0 *1 2.35,2.99
X$35 69 70 71 4 72 3 257 258 cell_2rw
* cell instance $36 m0 *1 3.525,2.99
X$36 73 74 75 4 76 3 257 258 cell_2rw
* cell instance $37 m0 *1 4.7,2.99
X$37 77 78 79 4 80 3 257 258 cell_2rw
* cell instance $38 m0 *1 5.875,2.99
X$38 81 82 83 4 84 3 257 258 cell_2rw
* cell instance $39 m0 *1 7.05,2.99
X$39 85 86 87 4 88 3 257 258 cell_2rw
* cell instance $40 m0 *1 8.225,2.99
X$40 89 90 91 4 92 3 257 258 cell_2rw
* cell instance $41 m0 *1 9.4,2.99
X$41 93 94 95 4 96 3 257 258 cell_2rw
* cell instance $42 m0 *1 10.575,2.99
X$42 97 98 99 4 100 3 257 258 cell_2rw
* cell instance $43 m0 *1 11.75,2.99
X$43 101 102 103 4 104 3 257 258 cell_2rw
* cell instance $44 m0 *1 12.925,2.99
X$44 105 106 107 4 108 3 257 258 cell_2rw
* cell instance $45 m0 *1 14.1,2.99
X$45 109 110 111 4 112 3 257 258 cell_2rw
* cell instance $46 m0 *1 15.275,2.99
X$46 113 114 115 4 116 3 257 258 cell_2rw
* cell instance $47 m0 *1 16.45,2.99
X$47 117 118 119 4 120 3 257 258 cell_2rw
* cell instance $48 m0 *1 17.625,2.99
X$48 121 122 123 4 124 3 257 258 cell_2rw
* cell instance $49 m0 *1 18.8,2.99
X$49 129 130 131 4 132 3 257 258 cell_2rw
* cell instance $50 m0 *1 19.975,2.99
X$50 133 134 135 4 136 3 257 258 cell_2rw
* cell instance $51 m0 *1 21.15,2.99
X$51 137 138 139 4 140 3 257 258 cell_2rw
* cell instance $52 m0 *1 22.325,2.99
X$52 141 142 143 4 144 3 257 258 cell_2rw
* cell instance $53 m0 *1 23.5,2.99
X$53 145 146 147 4 148 3 257 258 cell_2rw
* cell instance $54 m0 *1 24.675,2.99
X$54 149 150 151 4 152 3 257 258 cell_2rw
* cell instance $55 m0 *1 25.85,2.99
X$55 153 154 155 4 156 3 257 258 cell_2rw
* cell instance $56 m0 *1 27.025,2.99
X$56 157 158 159 4 160 3 257 258 cell_2rw
* cell instance $57 m0 *1 28.2,2.99
X$57 161 162 163 4 164 3 257 258 cell_2rw
* cell instance $58 m0 *1 29.375,2.99
X$58 165 166 167 4 168 3 257 258 cell_2rw
* cell instance $59 m0 *1 30.55,2.99
X$59 169 170 171 4 172 3 257 258 cell_2rw
* cell instance $60 m0 *1 31.725,2.99
X$60 173 174 175 4 176 3 257 258 cell_2rw
* cell instance $61 m0 *1 32.9,2.99
X$61 177 178 179 4 180 3 257 258 cell_2rw
* cell instance $62 m0 *1 34.075,2.99
X$62 181 182 183 4 184 3 257 258 cell_2rw
* cell instance $63 m0 *1 35.25,2.99
X$63 185 186 187 4 188 3 257 258 cell_2rw
* cell instance $64 m0 *1 36.425,2.99
X$64 189 190 191 4 192 3 257 258 cell_2rw
* cell instance $65 r0 *1 1.175,0
X$65 65 66 67 6 68 5 257 258 cell_2rw
* cell instance $66 r0 *1 0,0
X$66 61 62 63 6 64 5 257 258 cell_2rw
* cell instance $67 r0 *1 2.35,0
X$67 69 70 71 6 72 5 257 258 cell_2rw
* cell instance $68 r0 *1 3.525,0
X$68 73 74 75 6 76 5 257 258 cell_2rw
* cell instance $69 r0 *1 4.7,0
X$69 77 78 79 6 80 5 257 258 cell_2rw
* cell instance $70 r0 *1 5.875,0
X$70 81 82 83 6 84 5 257 258 cell_2rw
* cell instance $71 r0 *1 7.05,0
X$71 85 86 87 6 88 5 257 258 cell_2rw
* cell instance $72 r0 *1 8.225,0
X$72 89 90 91 6 92 5 257 258 cell_2rw
* cell instance $73 r0 *1 9.4,0
X$73 93 94 95 6 96 5 257 258 cell_2rw
* cell instance $74 r0 *1 10.575,0
X$74 97 98 99 6 100 5 257 258 cell_2rw
* cell instance $75 r0 *1 11.75,0
X$75 101 102 103 6 104 5 257 258 cell_2rw
* cell instance $76 r0 *1 12.925,0
X$76 105 106 107 6 108 5 257 258 cell_2rw
* cell instance $77 r0 *1 14.1,0
X$77 109 110 111 6 112 5 257 258 cell_2rw
* cell instance $78 r0 *1 15.275,0
X$78 113 114 115 6 116 5 257 258 cell_2rw
* cell instance $79 r0 *1 16.45,0
X$79 117 118 119 6 120 5 257 258 cell_2rw
* cell instance $80 r0 *1 17.625,0
X$80 121 122 123 6 124 5 257 258 cell_2rw
* cell instance $81 r0 *1 18.8,0
X$81 129 130 131 6 132 5 257 258 cell_2rw
* cell instance $82 r0 *1 19.975,0
X$82 133 134 135 6 136 5 257 258 cell_2rw
* cell instance $83 r0 *1 21.15,0
X$83 137 138 139 6 140 5 257 258 cell_2rw
* cell instance $84 r0 *1 22.325,0
X$84 141 142 143 6 144 5 257 258 cell_2rw
* cell instance $85 r0 *1 23.5,0
X$85 145 146 147 6 148 5 257 258 cell_2rw
* cell instance $86 r0 *1 24.675,0
X$86 149 150 151 6 152 5 257 258 cell_2rw
* cell instance $87 r0 *1 25.85,0
X$87 153 154 155 6 156 5 257 258 cell_2rw
* cell instance $88 r0 *1 27.025,0
X$88 157 158 159 6 160 5 257 258 cell_2rw
* cell instance $89 r0 *1 28.2,0
X$89 161 162 163 6 164 5 257 258 cell_2rw
* cell instance $90 r0 *1 29.375,0
X$90 165 166 167 6 168 5 257 258 cell_2rw
* cell instance $91 r0 *1 30.55,0
X$91 169 170 171 6 172 5 257 258 cell_2rw
* cell instance $92 r0 *1 31.725,0
X$92 173 174 175 6 176 5 257 258 cell_2rw
* cell instance $93 r0 *1 32.9,0
X$93 177 178 179 6 180 5 257 258 cell_2rw
* cell instance $94 r0 *1 34.075,0
X$94 181 182 183 6 184 5 257 258 cell_2rw
* cell instance $95 r0 *1 35.25,0
X$95 185 186 187 6 188 5 257 258 cell_2rw
* cell instance $96 r0 *1 36.425,0
X$96 189 190 191 6 192 5 257 258 cell_2rw
* cell instance $97 r0 *1 1.175,5.98
X$97 65 66 67 7 68 10 257 258 cell_2rw
* cell instance $98 r0 *1 0,5.98
X$98 61 62 63 7 64 10 257 258 cell_2rw
* cell instance $99 r0 *1 2.35,5.98
X$99 69 70 71 7 72 10 257 258 cell_2rw
* cell instance $100 r0 *1 3.525,5.98
X$100 73 74 75 7 76 10 257 258 cell_2rw
* cell instance $101 r0 *1 4.7,5.98
X$101 77 78 79 7 80 10 257 258 cell_2rw
* cell instance $102 r0 *1 5.875,5.98
X$102 81 82 83 7 84 10 257 258 cell_2rw
* cell instance $103 r0 *1 7.05,5.98
X$103 85 86 87 7 88 10 257 258 cell_2rw
* cell instance $104 r0 *1 8.225,5.98
X$104 89 90 91 7 92 10 257 258 cell_2rw
* cell instance $105 r0 *1 9.4,5.98
X$105 93 94 95 7 96 10 257 258 cell_2rw
* cell instance $106 r0 *1 10.575,5.98
X$106 97 98 99 7 100 10 257 258 cell_2rw
* cell instance $107 r0 *1 11.75,5.98
X$107 101 102 103 7 104 10 257 258 cell_2rw
* cell instance $108 r0 *1 12.925,5.98
X$108 105 106 107 7 108 10 257 258 cell_2rw
* cell instance $109 r0 *1 14.1,5.98
X$109 109 110 111 7 112 10 257 258 cell_2rw
* cell instance $110 r0 *1 15.275,5.98
X$110 113 114 115 7 116 10 257 258 cell_2rw
* cell instance $111 r0 *1 16.45,5.98
X$111 117 118 119 7 120 10 257 258 cell_2rw
* cell instance $112 r0 *1 17.625,5.98
X$112 121 122 123 7 124 10 257 258 cell_2rw
* cell instance $113 r0 *1 18.8,5.98
X$113 129 130 131 7 132 10 257 258 cell_2rw
* cell instance $114 r0 *1 19.975,5.98
X$114 133 134 135 7 136 10 257 258 cell_2rw
* cell instance $115 r0 *1 21.15,5.98
X$115 137 138 139 7 140 10 257 258 cell_2rw
* cell instance $116 r0 *1 22.325,5.98
X$116 141 142 143 7 144 10 257 258 cell_2rw
* cell instance $117 r0 *1 23.5,5.98
X$117 145 146 147 7 148 10 257 258 cell_2rw
* cell instance $118 r0 *1 24.675,5.98
X$118 149 150 151 7 152 10 257 258 cell_2rw
* cell instance $119 r0 *1 25.85,5.98
X$119 153 154 155 7 156 10 257 258 cell_2rw
* cell instance $120 r0 *1 27.025,5.98
X$120 157 158 159 7 160 10 257 258 cell_2rw
* cell instance $121 r0 *1 28.2,5.98
X$121 161 162 163 7 164 10 257 258 cell_2rw
* cell instance $122 r0 *1 29.375,5.98
X$122 165 166 167 7 168 10 257 258 cell_2rw
* cell instance $123 r0 *1 30.55,5.98
X$123 169 170 171 7 172 10 257 258 cell_2rw
* cell instance $124 r0 *1 31.725,5.98
X$124 173 174 175 7 176 10 257 258 cell_2rw
* cell instance $125 r0 *1 32.9,5.98
X$125 177 178 179 7 180 10 257 258 cell_2rw
* cell instance $126 r0 *1 34.075,5.98
X$126 181 182 183 7 184 10 257 258 cell_2rw
* cell instance $127 r0 *1 35.25,5.98
X$127 185 186 187 7 188 10 257 258 cell_2rw
* cell instance $128 r0 *1 36.425,5.98
X$128 189 190 191 7 192 10 257 258 cell_2rw
* cell instance $129 m0 *1 1.175,8.97
X$129 65 66 67 9 68 8 257 258 cell_2rw
* cell instance $130 m0 *1 0,8.97
X$130 61 62 63 9 64 8 257 258 cell_2rw
* cell instance $131 m0 *1 2.35,8.97
X$131 69 70 71 9 72 8 257 258 cell_2rw
* cell instance $132 m0 *1 3.525,8.97
X$132 73 74 75 9 76 8 257 258 cell_2rw
* cell instance $133 m0 *1 4.7,8.97
X$133 77 78 79 9 80 8 257 258 cell_2rw
* cell instance $134 m0 *1 5.875,8.97
X$134 81 82 83 9 84 8 257 258 cell_2rw
* cell instance $135 m0 *1 7.05,8.97
X$135 85 86 87 9 88 8 257 258 cell_2rw
* cell instance $136 m0 *1 8.225,8.97
X$136 89 90 91 9 92 8 257 258 cell_2rw
* cell instance $137 m0 *1 9.4,8.97
X$137 93 94 95 9 96 8 257 258 cell_2rw
* cell instance $138 m0 *1 10.575,8.97
X$138 97 98 99 9 100 8 257 258 cell_2rw
* cell instance $139 m0 *1 11.75,8.97
X$139 101 102 103 9 104 8 257 258 cell_2rw
* cell instance $140 m0 *1 12.925,8.97
X$140 105 106 107 9 108 8 257 258 cell_2rw
* cell instance $141 m0 *1 14.1,8.97
X$141 109 110 111 9 112 8 257 258 cell_2rw
* cell instance $142 m0 *1 15.275,8.97
X$142 113 114 115 9 116 8 257 258 cell_2rw
* cell instance $143 m0 *1 16.45,8.97
X$143 117 118 119 9 120 8 257 258 cell_2rw
* cell instance $144 m0 *1 17.625,8.97
X$144 121 122 123 9 124 8 257 258 cell_2rw
* cell instance $145 m0 *1 18.8,8.97
X$145 129 130 131 9 132 8 257 258 cell_2rw
* cell instance $146 m0 *1 19.975,8.97
X$146 133 134 135 9 136 8 257 258 cell_2rw
* cell instance $147 m0 *1 21.15,8.97
X$147 137 138 139 9 140 8 257 258 cell_2rw
* cell instance $148 m0 *1 22.325,8.97
X$148 141 142 143 9 144 8 257 258 cell_2rw
* cell instance $149 m0 *1 23.5,8.97
X$149 145 146 147 9 148 8 257 258 cell_2rw
* cell instance $150 m0 *1 24.675,8.97
X$150 149 150 151 9 152 8 257 258 cell_2rw
* cell instance $151 m0 *1 25.85,8.97
X$151 153 154 155 9 156 8 257 258 cell_2rw
* cell instance $152 m0 *1 27.025,8.97
X$152 157 158 159 9 160 8 257 258 cell_2rw
* cell instance $153 m0 *1 28.2,8.97
X$153 161 162 163 9 164 8 257 258 cell_2rw
* cell instance $154 m0 *1 29.375,8.97
X$154 165 166 167 9 168 8 257 258 cell_2rw
* cell instance $155 m0 *1 30.55,8.97
X$155 169 170 171 9 172 8 257 258 cell_2rw
* cell instance $156 m0 *1 31.725,8.97
X$156 173 174 175 9 176 8 257 258 cell_2rw
* cell instance $157 m0 *1 32.9,8.97
X$157 177 178 179 9 180 8 257 258 cell_2rw
* cell instance $158 m0 *1 34.075,8.97
X$158 181 182 183 9 184 8 257 258 cell_2rw
* cell instance $159 m0 *1 35.25,8.97
X$159 185 186 187 9 188 8 257 258 cell_2rw
* cell instance $160 m0 *1 36.425,8.97
X$160 189 190 191 9 192 8 257 258 cell_2rw
* cell instance $161 m0 *1 1.175,5.98
X$161 65 66 67 11 68 12 257 258 cell_2rw
* cell instance $162 m0 *1 0,5.98
X$162 61 62 63 11 64 12 257 258 cell_2rw
* cell instance $163 m0 *1 2.35,5.98
X$163 69 70 71 11 72 12 257 258 cell_2rw
* cell instance $164 m0 *1 3.525,5.98
X$164 73 74 75 11 76 12 257 258 cell_2rw
* cell instance $165 m0 *1 4.7,5.98
X$165 77 78 79 11 80 12 257 258 cell_2rw
* cell instance $166 m0 *1 5.875,5.98
X$166 81 82 83 11 84 12 257 258 cell_2rw
* cell instance $167 m0 *1 7.05,5.98
X$167 85 86 87 11 88 12 257 258 cell_2rw
* cell instance $168 m0 *1 8.225,5.98
X$168 89 90 91 11 92 12 257 258 cell_2rw
* cell instance $169 m0 *1 9.4,5.98
X$169 93 94 95 11 96 12 257 258 cell_2rw
* cell instance $170 m0 *1 10.575,5.98
X$170 97 98 99 11 100 12 257 258 cell_2rw
* cell instance $171 m0 *1 11.75,5.98
X$171 101 102 103 11 104 12 257 258 cell_2rw
* cell instance $172 m0 *1 12.925,5.98
X$172 105 106 107 11 108 12 257 258 cell_2rw
* cell instance $173 m0 *1 14.1,5.98
X$173 109 110 111 11 112 12 257 258 cell_2rw
* cell instance $174 m0 *1 15.275,5.98
X$174 113 114 115 11 116 12 257 258 cell_2rw
* cell instance $175 m0 *1 16.45,5.98
X$175 117 118 119 11 120 12 257 258 cell_2rw
* cell instance $176 m0 *1 17.625,5.98
X$176 121 122 123 11 124 12 257 258 cell_2rw
* cell instance $177 m0 *1 18.8,5.98
X$177 129 130 131 11 132 12 257 258 cell_2rw
* cell instance $178 m0 *1 19.975,5.98
X$178 133 134 135 11 136 12 257 258 cell_2rw
* cell instance $179 m0 *1 21.15,5.98
X$179 137 138 139 11 140 12 257 258 cell_2rw
* cell instance $180 m0 *1 22.325,5.98
X$180 141 142 143 11 144 12 257 258 cell_2rw
* cell instance $181 m0 *1 23.5,5.98
X$181 145 146 147 11 148 12 257 258 cell_2rw
* cell instance $182 m0 *1 24.675,5.98
X$182 149 150 151 11 152 12 257 258 cell_2rw
* cell instance $183 m0 *1 25.85,5.98
X$183 153 154 155 11 156 12 257 258 cell_2rw
* cell instance $184 m0 *1 27.025,5.98
X$184 157 158 159 11 160 12 257 258 cell_2rw
* cell instance $185 m0 *1 28.2,5.98
X$185 161 162 163 11 164 12 257 258 cell_2rw
* cell instance $186 m0 *1 29.375,5.98
X$186 165 166 167 11 168 12 257 258 cell_2rw
* cell instance $187 m0 *1 30.55,5.98
X$187 169 170 171 11 172 12 257 258 cell_2rw
* cell instance $188 m0 *1 31.725,5.98
X$188 173 174 175 11 176 12 257 258 cell_2rw
* cell instance $189 m0 *1 32.9,5.98
X$189 177 178 179 11 180 12 257 258 cell_2rw
* cell instance $190 m0 *1 34.075,5.98
X$190 181 182 183 11 184 12 257 258 cell_2rw
* cell instance $191 m0 *1 35.25,5.98
X$191 185 186 187 11 188 12 257 258 cell_2rw
* cell instance $192 m0 *1 36.425,5.98
X$192 189 190 191 11 192 12 257 258 cell_2rw
* cell instance $193 m0 *1 1.175,11.96
X$193 65 66 67 13 68 14 257 258 cell_2rw
* cell instance $194 m0 *1 0,11.96
X$194 61 62 63 13 64 14 257 258 cell_2rw
* cell instance $195 m0 *1 2.35,11.96
X$195 69 70 71 13 72 14 257 258 cell_2rw
* cell instance $196 m0 *1 3.525,11.96
X$196 73 74 75 13 76 14 257 258 cell_2rw
* cell instance $197 m0 *1 4.7,11.96
X$197 77 78 79 13 80 14 257 258 cell_2rw
* cell instance $198 m0 *1 5.875,11.96
X$198 81 82 83 13 84 14 257 258 cell_2rw
* cell instance $199 m0 *1 7.05,11.96
X$199 85 86 87 13 88 14 257 258 cell_2rw
* cell instance $200 m0 *1 8.225,11.96
X$200 89 90 91 13 92 14 257 258 cell_2rw
* cell instance $201 m0 *1 9.4,11.96
X$201 93 94 95 13 96 14 257 258 cell_2rw
* cell instance $202 m0 *1 10.575,11.96
X$202 97 98 99 13 100 14 257 258 cell_2rw
* cell instance $203 m0 *1 11.75,11.96
X$203 101 102 103 13 104 14 257 258 cell_2rw
* cell instance $204 m0 *1 12.925,11.96
X$204 105 106 107 13 108 14 257 258 cell_2rw
* cell instance $205 m0 *1 14.1,11.96
X$205 109 110 111 13 112 14 257 258 cell_2rw
* cell instance $206 m0 *1 15.275,11.96
X$206 113 114 115 13 116 14 257 258 cell_2rw
* cell instance $207 m0 *1 16.45,11.96
X$207 117 118 119 13 120 14 257 258 cell_2rw
* cell instance $208 m0 *1 17.625,11.96
X$208 121 122 123 13 124 14 257 258 cell_2rw
* cell instance $209 m0 *1 18.8,11.96
X$209 129 130 131 13 132 14 257 258 cell_2rw
* cell instance $210 m0 *1 19.975,11.96
X$210 133 134 135 13 136 14 257 258 cell_2rw
* cell instance $211 m0 *1 21.15,11.96
X$211 137 138 139 13 140 14 257 258 cell_2rw
* cell instance $212 m0 *1 22.325,11.96
X$212 141 142 143 13 144 14 257 258 cell_2rw
* cell instance $213 m0 *1 23.5,11.96
X$213 145 146 147 13 148 14 257 258 cell_2rw
* cell instance $214 m0 *1 24.675,11.96
X$214 149 150 151 13 152 14 257 258 cell_2rw
* cell instance $215 m0 *1 25.85,11.96
X$215 153 154 155 13 156 14 257 258 cell_2rw
* cell instance $216 m0 *1 27.025,11.96
X$216 157 158 159 13 160 14 257 258 cell_2rw
* cell instance $217 m0 *1 28.2,11.96
X$217 161 162 163 13 164 14 257 258 cell_2rw
* cell instance $218 m0 *1 29.375,11.96
X$218 165 166 167 13 168 14 257 258 cell_2rw
* cell instance $219 m0 *1 30.55,11.96
X$219 169 170 171 13 172 14 257 258 cell_2rw
* cell instance $220 m0 *1 31.725,11.96
X$220 173 174 175 13 176 14 257 258 cell_2rw
* cell instance $221 m0 *1 32.9,11.96
X$221 177 178 179 13 180 14 257 258 cell_2rw
* cell instance $222 m0 *1 34.075,11.96
X$222 181 182 183 13 184 14 257 258 cell_2rw
* cell instance $223 m0 *1 35.25,11.96
X$223 185 186 187 13 188 14 257 258 cell_2rw
* cell instance $224 m0 *1 36.425,11.96
X$224 189 190 191 13 192 14 257 258 cell_2rw
* cell instance $225 r0 *1 1.175,11.96
X$225 65 66 67 16 68 15 257 258 cell_2rw
* cell instance $226 r0 *1 0,11.96
X$226 61 62 63 16 64 15 257 258 cell_2rw
* cell instance $227 r0 *1 2.35,11.96
X$227 69 70 71 16 72 15 257 258 cell_2rw
* cell instance $228 r0 *1 3.525,11.96
X$228 73 74 75 16 76 15 257 258 cell_2rw
* cell instance $229 r0 *1 4.7,11.96
X$229 77 78 79 16 80 15 257 258 cell_2rw
* cell instance $230 r0 *1 5.875,11.96
X$230 81 82 83 16 84 15 257 258 cell_2rw
* cell instance $231 r0 *1 7.05,11.96
X$231 85 86 87 16 88 15 257 258 cell_2rw
* cell instance $232 r0 *1 8.225,11.96
X$232 89 90 91 16 92 15 257 258 cell_2rw
* cell instance $233 r0 *1 9.4,11.96
X$233 93 94 95 16 96 15 257 258 cell_2rw
* cell instance $234 r0 *1 10.575,11.96
X$234 97 98 99 16 100 15 257 258 cell_2rw
* cell instance $235 r0 *1 11.75,11.96
X$235 101 102 103 16 104 15 257 258 cell_2rw
* cell instance $236 r0 *1 12.925,11.96
X$236 105 106 107 16 108 15 257 258 cell_2rw
* cell instance $237 r0 *1 14.1,11.96
X$237 109 110 111 16 112 15 257 258 cell_2rw
* cell instance $238 r0 *1 15.275,11.96
X$238 113 114 115 16 116 15 257 258 cell_2rw
* cell instance $239 r0 *1 16.45,11.96
X$239 117 118 119 16 120 15 257 258 cell_2rw
* cell instance $240 r0 *1 17.625,11.96
X$240 121 122 123 16 124 15 257 258 cell_2rw
* cell instance $241 r0 *1 18.8,11.96
X$241 129 130 131 16 132 15 257 258 cell_2rw
* cell instance $242 r0 *1 19.975,11.96
X$242 133 134 135 16 136 15 257 258 cell_2rw
* cell instance $243 r0 *1 21.15,11.96
X$243 137 138 139 16 140 15 257 258 cell_2rw
* cell instance $244 r0 *1 22.325,11.96
X$244 141 142 143 16 144 15 257 258 cell_2rw
* cell instance $245 r0 *1 23.5,11.96
X$245 145 146 147 16 148 15 257 258 cell_2rw
* cell instance $246 r0 *1 24.675,11.96
X$246 149 150 151 16 152 15 257 258 cell_2rw
* cell instance $247 r0 *1 25.85,11.96
X$247 153 154 155 16 156 15 257 258 cell_2rw
* cell instance $248 r0 *1 27.025,11.96
X$248 157 158 159 16 160 15 257 258 cell_2rw
* cell instance $249 r0 *1 28.2,11.96
X$249 161 162 163 16 164 15 257 258 cell_2rw
* cell instance $250 r0 *1 29.375,11.96
X$250 165 166 167 16 168 15 257 258 cell_2rw
* cell instance $251 r0 *1 30.55,11.96
X$251 169 170 171 16 172 15 257 258 cell_2rw
* cell instance $252 r0 *1 31.725,11.96
X$252 173 174 175 16 176 15 257 258 cell_2rw
* cell instance $253 r0 *1 32.9,11.96
X$253 177 178 179 16 180 15 257 258 cell_2rw
* cell instance $254 r0 *1 34.075,11.96
X$254 181 182 183 16 184 15 257 258 cell_2rw
* cell instance $255 r0 *1 35.25,11.96
X$255 185 186 187 16 188 15 257 258 cell_2rw
* cell instance $256 r0 *1 36.425,11.96
X$256 189 190 191 16 192 15 257 258 cell_2rw
* cell instance $257 r0 *1 1.175,8.97
X$257 65 66 67 17 68 18 257 258 cell_2rw
* cell instance $258 r0 *1 0,8.97
X$258 61 62 63 17 64 18 257 258 cell_2rw
* cell instance $259 r0 *1 2.35,8.97
X$259 69 70 71 17 72 18 257 258 cell_2rw
* cell instance $260 r0 *1 3.525,8.97
X$260 73 74 75 17 76 18 257 258 cell_2rw
* cell instance $261 r0 *1 4.7,8.97
X$261 77 78 79 17 80 18 257 258 cell_2rw
* cell instance $262 r0 *1 5.875,8.97
X$262 81 82 83 17 84 18 257 258 cell_2rw
* cell instance $263 r0 *1 7.05,8.97
X$263 85 86 87 17 88 18 257 258 cell_2rw
* cell instance $264 r0 *1 8.225,8.97
X$264 89 90 91 17 92 18 257 258 cell_2rw
* cell instance $265 r0 *1 9.4,8.97
X$265 93 94 95 17 96 18 257 258 cell_2rw
* cell instance $266 r0 *1 10.575,8.97
X$266 97 98 99 17 100 18 257 258 cell_2rw
* cell instance $267 r0 *1 11.75,8.97
X$267 101 102 103 17 104 18 257 258 cell_2rw
* cell instance $268 r0 *1 12.925,8.97
X$268 105 106 107 17 108 18 257 258 cell_2rw
* cell instance $269 r0 *1 14.1,8.97
X$269 109 110 111 17 112 18 257 258 cell_2rw
* cell instance $270 r0 *1 15.275,8.97
X$270 113 114 115 17 116 18 257 258 cell_2rw
* cell instance $271 r0 *1 16.45,8.97
X$271 117 118 119 17 120 18 257 258 cell_2rw
* cell instance $272 r0 *1 17.625,8.97
X$272 121 122 123 17 124 18 257 258 cell_2rw
* cell instance $273 r0 *1 18.8,8.97
X$273 129 130 131 17 132 18 257 258 cell_2rw
* cell instance $274 r0 *1 19.975,8.97
X$274 133 134 135 17 136 18 257 258 cell_2rw
* cell instance $275 r0 *1 21.15,8.97
X$275 137 138 139 17 140 18 257 258 cell_2rw
* cell instance $276 r0 *1 22.325,8.97
X$276 141 142 143 17 144 18 257 258 cell_2rw
* cell instance $277 r0 *1 23.5,8.97
X$277 145 146 147 17 148 18 257 258 cell_2rw
* cell instance $278 r0 *1 24.675,8.97
X$278 149 150 151 17 152 18 257 258 cell_2rw
* cell instance $279 r0 *1 25.85,8.97
X$279 153 154 155 17 156 18 257 258 cell_2rw
* cell instance $280 r0 *1 27.025,8.97
X$280 157 158 159 17 160 18 257 258 cell_2rw
* cell instance $281 r0 *1 28.2,8.97
X$281 161 162 163 17 164 18 257 258 cell_2rw
* cell instance $282 r0 *1 29.375,8.97
X$282 165 166 167 17 168 18 257 258 cell_2rw
* cell instance $283 r0 *1 30.55,8.97
X$283 169 170 171 17 172 18 257 258 cell_2rw
* cell instance $284 r0 *1 31.725,8.97
X$284 173 174 175 17 176 18 257 258 cell_2rw
* cell instance $285 r0 *1 32.9,8.97
X$285 177 178 179 17 180 18 257 258 cell_2rw
* cell instance $286 r0 *1 34.075,8.97
X$286 181 182 183 17 184 18 257 258 cell_2rw
* cell instance $287 r0 *1 35.25,8.97
X$287 185 186 187 17 188 18 257 258 cell_2rw
* cell instance $288 r0 *1 36.425,8.97
X$288 189 190 191 17 192 18 257 258 cell_2rw
* cell instance $289 r0 *1 1.175,14.95
X$289 65 66 67 20 68 19 257 258 cell_2rw
* cell instance $290 r0 *1 0,14.95
X$290 61 62 63 20 64 19 257 258 cell_2rw
* cell instance $291 r0 *1 2.35,14.95
X$291 69 70 71 20 72 19 257 258 cell_2rw
* cell instance $292 r0 *1 3.525,14.95
X$292 73 74 75 20 76 19 257 258 cell_2rw
* cell instance $293 r0 *1 4.7,14.95
X$293 77 78 79 20 80 19 257 258 cell_2rw
* cell instance $294 r0 *1 5.875,14.95
X$294 81 82 83 20 84 19 257 258 cell_2rw
* cell instance $295 r0 *1 7.05,14.95
X$295 85 86 87 20 88 19 257 258 cell_2rw
* cell instance $296 r0 *1 8.225,14.95
X$296 89 90 91 20 92 19 257 258 cell_2rw
* cell instance $297 r0 *1 9.4,14.95
X$297 93 94 95 20 96 19 257 258 cell_2rw
* cell instance $298 r0 *1 10.575,14.95
X$298 97 98 99 20 100 19 257 258 cell_2rw
* cell instance $299 r0 *1 11.75,14.95
X$299 101 102 103 20 104 19 257 258 cell_2rw
* cell instance $300 r0 *1 12.925,14.95
X$300 105 106 107 20 108 19 257 258 cell_2rw
* cell instance $301 r0 *1 14.1,14.95
X$301 109 110 111 20 112 19 257 258 cell_2rw
* cell instance $302 r0 *1 15.275,14.95
X$302 113 114 115 20 116 19 257 258 cell_2rw
* cell instance $303 r0 *1 16.45,14.95
X$303 117 118 119 20 120 19 257 258 cell_2rw
* cell instance $304 r0 *1 17.625,14.95
X$304 121 122 123 20 124 19 257 258 cell_2rw
* cell instance $305 r0 *1 18.8,14.95
X$305 129 130 131 20 132 19 257 258 cell_2rw
* cell instance $306 r0 *1 19.975,14.95
X$306 133 134 135 20 136 19 257 258 cell_2rw
* cell instance $307 r0 *1 21.15,14.95
X$307 137 138 139 20 140 19 257 258 cell_2rw
* cell instance $308 r0 *1 22.325,14.95
X$308 141 142 143 20 144 19 257 258 cell_2rw
* cell instance $309 r0 *1 23.5,14.95
X$309 145 146 147 20 148 19 257 258 cell_2rw
* cell instance $310 r0 *1 24.675,14.95
X$310 149 150 151 20 152 19 257 258 cell_2rw
* cell instance $311 r0 *1 25.85,14.95
X$311 153 154 155 20 156 19 257 258 cell_2rw
* cell instance $312 r0 *1 27.025,14.95
X$312 157 158 159 20 160 19 257 258 cell_2rw
* cell instance $313 r0 *1 28.2,14.95
X$313 161 162 163 20 164 19 257 258 cell_2rw
* cell instance $314 r0 *1 29.375,14.95
X$314 165 166 167 20 168 19 257 258 cell_2rw
* cell instance $315 r0 *1 30.55,14.95
X$315 169 170 171 20 172 19 257 258 cell_2rw
* cell instance $316 r0 *1 31.725,14.95
X$316 173 174 175 20 176 19 257 258 cell_2rw
* cell instance $317 r0 *1 32.9,14.95
X$317 177 178 179 20 180 19 257 258 cell_2rw
* cell instance $318 r0 *1 34.075,14.95
X$318 181 182 183 20 184 19 257 258 cell_2rw
* cell instance $319 r0 *1 35.25,14.95
X$319 185 186 187 20 188 19 257 258 cell_2rw
* cell instance $320 r0 *1 36.425,14.95
X$320 189 190 191 20 192 19 257 258 cell_2rw
* cell instance $321 m0 *1 1.175,17.94
X$321 65 66 67 21 68 22 257 258 cell_2rw
* cell instance $322 m0 *1 0,17.94
X$322 61 62 63 21 64 22 257 258 cell_2rw
* cell instance $323 m0 *1 2.35,17.94
X$323 69 70 71 21 72 22 257 258 cell_2rw
* cell instance $324 m0 *1 3.525,17.94
X$324 73 74 75 21 76 22 257 258 cell_2rw
* cell instance $325 m0 *1 4.7,17.94
X$325 77 78 79 21 80 22 257 258 cell_2rw
* cell instance $326 m0 *1 5.875,17.94
X$326 81 82 83 21 84 22 257 258 cell_2rw
* cell instance $327 m0 *1 7.05,17.94
X$327 85 86 87 21 88 22 257 258 cell_2rw
* cell instance $328 m0 *1 8.225,17.94
X$328 89 90 91 21 92 22 257 258 cell_2rw
* cell instance $329 m0 *1 9.4,17.94
X$329 93 94 95 21 96 22 257 258 cell_2rw
* cell instance $330 m0 *1 10.575,17.94
X$330 97 98 99 21 100 22 257 258 cell_2rw
* cell instance $331 m0 *1 11.75,17.94
X$331 101 102 103 21 104 22 257 258 cell_2rw
* cell instance $332 m0 *1 12.925,17.94
X$332 105 106 107 21 108 22 257 258 cell_2rw
* cell instance $333 m0 *1 14.1,17.94
X$333 109 110 111 21 112 22 257 258 cell_2rw
* cell instance $334 m0 *1 15.275,17.94
X$334 113 114 115 21 116 22 257 258 cell_2rw
* cell instance $335 m0 *1 16.45,17.94
X$335 117 118 119 21 120 22 257 258 cell_2rw
* cell instance $336 m0 *1 17.625,17.94
X$336 121 122 123 21 124 22 257 258 cell_2rw
* cell instance $337 m0 *1 18.8,17.94
X$337 129 130 131 21 132 22 257 258 cell_2rw
* cell instance $338 m0 *1 19.975,17.94
X$338 133 134 135 21 136 22 257 258 cell_2rw
* cell instance $339 m0 *1 21.15,17.94
X$339 137 138 139 21 140 22 257 258 cell_2rw
* cell instance $340 m0 *1 22.325,17.94
X$340 141 142 143 21 144 22 257 258 cell_2rw
* cell instance $341 m0 *1 23.5,17.94
X$341 145 146 147 21 148 22 257 258 cell_2rw
* cell instance $342 m0 *1 24.675,17.94
X$342 149 150 151 21 152 22 257 258 cell_2rw
* cell instance $343 m0 *1 25.85,17.94
X$343 153 154 155 21 156 22 257 258 cell_2rw
* cell instance $344 m0 *1 27.025,17.94
X$344 157 158 159 21 160 22 257 258 cell_2rw
* cell instance $345 m0 *1 28.2,17.94
X$345 161 162 163 21 164 22 257 258 cell_2rw
* cell instance $346 m0 *1 29.375,17.94
X$346 165 166 167 21 168 22 257 258 cell_2rw
* cell instance $347 m0 *1 30.55,17.94
X$347 169 170 171 21 172 22 257 258 cell_2rw
* cell instance $348 m0 *1 31.725,17.94
X$348 173 174 175 21 176 22 257 258 cell_2rw
* cell instance $349 m0 *1 32.9,17.94
X$349 177 178 179 21 180 22 257 258 cell_2rw
* cell instance $350 m0 *1 34.075,17.94
X$350 181 182 183 21 184 22 257 258 cell_2rw
* cell instance $351 m0 *1 35.25,17.94
X$351 185 186 187 21 188 22 257 258 cell_2rw
* cell instance $352 m0 *1 36.425,17.94
X$352 189 190 191 21 192 22 257 258 cell_2rw
* cell instance $353 m0 *1 1.175,14.95
X$353 65 66 67 24 68 23 257 258 cell_2rw
* cell instance $354 m0 *1 0,14.95
X$354 61 62 63 24 64 23 257 258 cell_2rw
* cell instance $355 m0 *1 2.35,14.95
X$355 69 70 71 24 72 23 257 258 cell_2rw
* cell instance $356 m0 *1 3.525,14.95
X$356 73 74 75 24 76 23 257 258 cell_2rw
* cell instance $357 m0 *1 4.7,14.95
X$357 77 78 79 24 80 23 257 258 cell_2rw
* cell instance $358 m0 *1 5.875,14.95
X$358 81 82 83 24 84 23 257 258 cell_2rw
* cell instance $359 m0 *1 7.05,14.95
X$359 85 86 87 24 88 23 257 258 cell_2rw
* cell instance $360 m0 *1 8.225,14.95
X$360 89 90 91 24 92 23 257 258 cell_2rw
* cell instance $361 m0 *1 9.4,14.95
X$361 93 94 95 24 96 23 257 258 cell_2rw
* cell instance $362 m0 *1 10.575,14.95
X$362 97 98 99 24 100 23 257 258 cell_2rw
* cell instance $363 m0 *1 11.75,14.95
X$363 101 102 103 24 104 23 257 258 cell_2rw
* cell instance $364 m0 *1 12.925,14.95
X$364 105 106 107 24 108 23 257 258 cell_2rw
* cell instance $365 m0 *1 14.1,14.95
X$365 109 110 111 24 112 23 257 258 cell_2rw
* cell instance $366 m0 *1 15.275,14.95
X$366 113 114 115 24 116 23 257 258 cell_2rw
* cell instance $367 m0 *1 16.45,14.95
X$367 117 118 119 24 120 23 257 258 cell_2rw
* cell instance $368 m0 *1 17.625,14.95
X$368 121 122 123 24 124 23 257 258 cell_2rw
* cell instance $369 m0 *1 18.8,14.95
X$369 129 130 131 24 132 23 257 258 cell_2rw
* cell instance $370 m0 *1 19.975,14.95
X$370 133 134 135 24 136 23 257 258 cell_2rw
* cell instance $371 m0 *1 21.15,14.95
X$371 137 138 139 24 140 23 257 258 cell_2rw
* cell instance $372 m0 *1 22.325,14.95
X$372 141 142 143 24 144 23 257 258 cell_2rw
* cell instance $373 m0 *1 23.5,14.95
X$373 145 146 147 24 148 23 257 258 cell_2rw
* cell instance $374 m0 *1 24.675,14.95
X$374 149 150 151 24 152 23 257 258 cell_2rw
* cell instance $375 m0 *1 25.85,14.95
X$375 153 154 155 24 156 23 257 258 cell_2rw
* cell instance $376 m0 *1 27.025,14.95
X$376 157 158 159 24 160 23 257 258 cell_2rw
* cell instance $377 m0 *1 28.2,14.95
X$377 161 162 163 24 164 23 257 258 cell_2rw
* cell instance $378 m0 *1 29.375,14.95
X$378 165 166 167 24 168 23 257 258 cell_2rw
* cell instance $379 m0 *1 30.55,14.95
X$379 169 170 171 24 172 23 257 258 cell_2rw
* cell instance $380 m0 *1 31.725,14.95
X$380 173 174 175 24 176 23 257 258 cell_2rw
* cell instance $381 m0 *1 32.9,14.95
X$381 177 178 179 24 180 23 257 258 cell_2rw
* cell instance $382 m0 *1 34.075,14.95
X$382 181 182 183 24 184 23 257 258 cell_2rw
* cell instance $383 m0 *1 35.25,14.95
X$383 185 186 187 24 188 23 257 258 cell_2rw
* cell instance $384 m0 *1 36.425,14.95
X$384 189 190 191 24 192 23 257 258 cell_2rw
* cell instance $385 r0 *1 1.175,20.93
X$385 65 66 67 28 68 25 257 258 cell_2rw
* cell instance $386 r0 *1 0,20.93
X$386 61 62 63 28 64 25 257 258 cell_2rw
* cell instance $387 r0 *1 2.35,20.93
X$387 69 70 71 28 72 25 257 258 cell_2rw
* cell instance $388 r0 *1 3.525,20.93
X$388 73 74 75 28 76 25 257 258 cell_2rw
* cell instance $389 r0 *1 4.7,20.93
X$389 77 78 79 28 80 25 257 258 cell_2rw
* cell instance $390 r0 *1 5.875,20.93
X$390 81 82 83 28 84 25 257 258 cell_2rw
* cell instance $391 r0 *1 7.05,20.93
X$391 85 86 87 28 88 25 257 258 cell_2rw
* cell instance $392 r0 *1 8.225,20.93
X$392 89 90 91 28 92 25 257 258 cell_2rw
* cell instance $393 r0 *1 9.4,20.93
X$393 93 94 95 28 96 25 257 258 cell_2rw
* cell instance $394 r0 *1 10.575,20.93
X$394 97 98 99 28 100 25 257 258 cell_2rw
* cell instance $395 r0 *1 11.75,20.93
X$395 101 102 103 28 104 25 257 258 cell_2rw
* cell instance $396 r0 *1 12.925,20.93
X$396 105 106 107 28 108 25 257 258 cell_2rw
* cell instance $397 r0 *1 14.1,20.93
X$397 109 110 111 28 112 25 257 258 cell_2rw
* cell instance $398 r0 *1 15.275,20.93
X$398 113 114 115 28 116 25 257 258 cell_2rw
* cell instance $399 r0 *1 16.45,20.93
X$399 117 118 119 28 120 25 257 258 cell_2rw
* cell instance $400 r0 *1 17.625,20.93
X$400 121 122 123 28 124 25 257 258 cell_2rw
* cell instance $401 r0 *1 18.8,20.93
X$401 129 130 131 28 132 25 257 258 cell_2rw
* cell instance $402 r0 *1 19.975,20.93
X$402 133 134 135 28 136 25 257 258 cell_2rw
* cell instance $403 r0 *1 21.15,20.93
X$403 137 138 139 28 140 25 257 258 cell_2rw
* cell instance $404 r0 *1 22.325,20.93
X$404 141 142 143 28 144 25 257 258 cell_2rw
* cell instance $405 r0 *1 23.5,20.93
X$405 145 146 147 28 148 25 257 258 cell_2rw
* cell instance $406 r0 *1 24.675,20.93
X$406 149 150 151 28 152 25 257 258 cell_2rw
* cell instance $407 r0 *1 25.85,20.93
X$407 153 154 155 28 156 25 257 258 cell_2rw
* cell instance $408 r0 *1 27.025,20.93
X$408 157 158 159 28 160 25 257 258 cell_2rw
* cell instance $409 r0 *1 28.2,20.93
X$409 161 162 163 28 164 25 257 258 cell_2rw
* cell instance $410 r0 *1 29.375,20.93
X$410 165 166 167 28 168 25 257 258 cell_2rw
* cell instance $411 r0 *1 30.55,20.93
X$411 169 170 171 28 172 25 257 258 cell_2rw
* cell instance $412 r0 *1 31.725,20.93
X$412 173 174 175 28 176 25 257 258 cell_2rw
* cell instance $413 r0 *1 32.9,20.93
X$413 177 178 179 28 180 25 257 258 cell_2rw
* cell instance $414 r0 *1 34.075,20.93
X$414 181 182 183 28 184 25 257 258 cell_2rw
* cell instance $415 r0 *1 35.25,20.93
X$415 185 186 187 28 188 25 257 258 cell_2rw
* cell instance $416 r0 *1 36.425,20.93
X$416 189 190 191 28 192 25 257 258 cell_2rw
* cell instance $417 m0 *1 1.175,20.93
X$417 65 66 67 26 68 29 257 258 cell_2rw
* cell instance $418 m0 *1 0,20.93
X$418 61 62 63 26 64 29 257 258 cell_2rw
* cell instance $419 m0 *1 2.35,20.93
X$419 69 70 71 26 72 29 257 258 cell_2rw
* cell instance $420 m0 *1 3.525,20.93
X$420 73 74 75 26 76 29 257 258 cell_2rw
* cell instance $421 m0 *1 4.7,20.93
X$421 77 78 79 26 80 29 257 258 cell_2rw
* cell instance $422 m0 *1 5.875,20.93
X$422 81 82 83 26 84 29 257 258 cell_2rw
* cell instance $423 m0 *1 7.05,20.93
X$423 85 86 87 26 88 29 257 258 cell_2rw
* cell instance $424 m0 *1 8.225,20.93
X$424 89 90 91 26 92 29 257 258 cell_2rw
* cell instance $425 m0 *1 9.4,20.93
X$425 93 94 95 26 96 29 257 258 cell_2rw
* cell instance $426 m0 *1 10.575,20.93
X$426 97 98 99 26 100 29 257 258 cell_2rw
* cell instance $427 m0 *1 11.75,20.93
X$427 101 102 103 26 104 29 257 258 cell_2rw
* cell instance $428 m0 *1 12.925,20.93
X$428 105 106 107 26 108 29 257 258 cell_2rw
* cell instance $429 m0 *1 14.1,20.93
X$429 109 110 111 26 112 29 257 258 cell_2rw
* cell instance $430 m0 *1 15.275,20.93
X$430 113 114 115 26 116 29 257 258 cell_2rw
* cell instance $431 m0 *1 16.45,20.93
X$431 117 118 119 26 120 29 257 258 cell_2rw
* cell instance $432 m0 *1 17.625,20.93
X$432 121 122 123 26 124 29 257 258 cell_2rw
* cell instance $433 m0 *1 18.8,20.93
X$433 129 130 131 26 132 29 257 258 cell_2rw
* cell instance $434 m0 *1 19.975,20.93
X$434 133 134 135 26 136 29 257 258 cell_2rw
* cell instance $435 m0 *1 21.15,20.93
X$435 137 138 139 26 140 29 257 258 cell_2rw
* cell instance $436 m0 *1 22.325,20.93
X$436 141 142 143 26 144 29 257 258 cell_2rw
* cell instance $437 m0 *1 23.5,20.93
X$437 145 146 147 26 148 29 257 258 cell_2rw
* cell instance $438 m0 *1 24.675,20.93
X$438 149 150 151 26 152 29 257 258 cell_2rw
* cell instance $439 m0 *1 25.85,20.93
X$439 153 154 155 26 156 29 257 258 cell_2rw
* cell instance $440 m0 *1 27.025,20.93
X$440 157 158 159 26 160 29 257 258 cell_2rw
* cell instance $441 m0 *1 28.2,20.93
X$441 161 162 163 26 164 29 257 258 cell_2rw
* cell instance $442 m0 *1 29.375,20.93
X$442 165 166 167 26 168 29 257 258 cell_2rw
* cell instance $443 m0 *1 30.55,20.93
X$443 169 170 171 26 172 29 257 258 cell_2rw
* cell instance $444 m0 *1 31.725,20.93
X$444 173 174 175 26 176 29 257 258 cell_2rw
* cell instance $445 m0 *1 32.9,20.93
X$445 177 178 179 26 180 29 257 258 cell_2rw
* cell instance $446 m0 *1 34.075,20.93
X$446 181 182 183 26 184 29 257 258 cell_2rw
* cell instance $447 m0 *1 35.25,20.93
X$447 185 186 187 26 188 29 257 258 cell_2rw
* cell instance $448 m0 *1 36.425,20.93
X$448 189 190 191 26 192 29 257 258 cell_2rw
* cell instance $449 r0 *1 1.175,17.94
X$449 65 66 67 27 68 30 257 258 cell_2rw
* cell instance $450 r0 *1 0,17.94
X$450 61 62 63 27 64 30 257 258 cell_2rw
* cell instance $451 r0 *1 2.35,17.94
X$451 69 70 71 27 72 30 257 258 cell_2rw
* cell instance $452 r0 *1 3.525,17.94
X$452 73 74 75 27 76 30 257 258 cell_2rw
* cell instance $453 r0 *1 4.7,17.94
X$453 77 78 79 27 80 30 257 258 cell_2rw
* cell instance $454 r0 *1 5.875,17.94
X$454 81 82 83 27 84 30 257 258 cell_2rw
* cell instance $455 r0 *1 7.05,17.94
X$455 85 86 87 27 88 30 257 258 cell_2rw
* cell instance $456 r0 *1 8.225,17.94
X$456 89 90 91 27 92 30 257 258 cell_2rw
* cell instance $457 r0 *1 9.4,17.94
X$457 93 94 95 27 96 30 257 258 cell_2rw
* cell instance $458 r0 *1 10.575,17.94
X$458 97 98 99 27 100 30 257 258 cell_2rw
* cell instance $459 r0 *1 11.75,17.94
X$459 101 102 103 27 104 30 257 258 cell_2rw
* cell instance $460 r0 *1 12.925,17.94
X$460 105 106 107 27 108 30 257 258 cell_2rw
* cell instance $461 r0 *1 14.1,17.94
X$461 109 110 111 27 112 30 257 258 cell_2rw
* cell instance $462 r0 *1 15.275,17.94
X$462 113 114 115 27 116 30 257 258 cell_2rw
* cell instance $463 r0 *1 16.45,17.94
X$463 117 118 119 27 120 30 257 258 cell_2rw
* cell instance $464 r0 *1 17.625,17.94
X$464 121 122 123 27 124 30 257 258 cell_2rw
* cell instance $465 r0 *1 18.8,17.94
X$465 129 130 131 27 132 30 257 258 cell_2rw
* cell instance $466 r0 *1 19.975,17.94
X$466 133 134 135 27 136 30 257 258 cell_2rw
* cell instance $467 r0 *1 21.15,17.94
X$467 137 138 139 27 140 30 257 258 cell_2rw
* cell instance $468 r0 *1 22.325,17.94
X$468 141 142 143 27 144 30 257 258 cell_2rw
* cell instance $469 r0 *1 23.5,17.94
X$469 145 146 147 27 148 30 257 258 cell_2rw
* cell instance $470 r0 *1 24.675,17.94
X$470 149 150 151 27 152 30 257 258 cell_2rw
* cell instance $471 r0 *1 25.85,17.94
X$471 153 154 155 27 156 30 257 258 cell_2rw
* cell instance $472 r0 *1 27.025,17.94
X$472 157 158 159 27 160 30 257 258 cell_2rw
* cell instance $473 r0 *1 28.2,17.94
X$473 161 162 163 27 164 30 257 258 cell_2rw
* cell instance $474 r0 *1 29.375,17.94
X$474 165 166 167 27 168 30 257 258 cell_2rw
* cell instance $475 r0 *1 30.55,17.94
X$475 169 170 171 27 172 30 257 258 cell_2rw
* cell instance $476 r0 *1 31.725,17.94
X$476 173 174 175 27 176 30 257 258 cell_2rw
* cell instance $477 r0 *1 32.9,17.94
X$477 177 178 179 27 180 30 257 258 cell_2rw
* cell instance $478 r0 *1 34.075,17.94
X$478 181 182 183 27 184 30 257 258 cell_2rw
* cell instance $479 r0 *1 35.25,17.94
X$479 185 186 187 27 188 30 257 258 cell_2rw
* cell instance $480 r0 *1 36.425,17.94
X$480 189 190 191 27 192 30 257 258 cell_2rw
* cell instance $481 r0 *1 1.175,23.92
X$481 65 66 67 31 68 33 257 258 cell_2rw
* cell instance $482 r0 *1 0,23.92
X$482 61 62 63 31 64 33 257 258 cell_2rw
* cell instance $483 r0 *1 2.35,23.92
X$483 69 70 71 31 72 33 257 258 cell_2rw
* cell instance $484 r0 *1 3.525,23.92
X$484 73 74 75 31 76 33 257 258 cell_2rw
* cell instance $485 r0 *1 4.7,23.92
X$485 77 78 79 31 80 33 257 258 cell_2rw
* cell instance $486 r0 *1 5.875,23.92
X$486 81 82 83 31 84 33 257 258 cell_2rw
* cell instance $487 r0 *1 7.05,23.92
X$487 85 86 87 31 88 33 257 258 cell_2rw
* cell instance $488 r0 *1 8.225,23.92
X$488 89 90 91 31 92 33 257 258 cell_2rw
* cell instance $489 r0 *1 9.4,23.92
X$489 93 94 95 31 96 33 257 258 cell_2rw
* cell instance $490 r0 *1 10.575,23.92
X$490 97 98 99 31 100 33 257 258 cell_2rw
* cell instance $491 r0 *1 11.75,23.92
X$491 101 102 103 31 104 33 257 258 cell_2rw
* cell instance $492 r0 *1 12.925,23.92
X$492 105 106 107 31 108 33 257 258 cell_2rw
* cell instance $493 r0 *1 14.1,23.92
X$493 109 110 111 31 112 33 257 258 cell_2rw
* cell instance $494 r0 *1 15.275,23.92
X$494 113 114 115 31 116 33 257 258 cell_2rw
* cell instance $495 r0 *1 16.45,23.92
X$495 117 118 119 31 120 33 257 258 cell_2rw
* cell instance $496 r0 *1 17.625,23.92
X$496 121 122 123 31 124 33 257 258 cell_2rw
* cell instance $497 r0 *1 18.8,23.92
X$497 129 130 131 31 132 33 257 258 cell_2rw
* cell instance $498 r0 *1 19.975,23.92
X$498 133 134 135 31 136 33 257 258 cell_2rw
* cell instance $499 r0 *1 21.15,23.92
X$499 137 138 139 31 140 33 257 258 cell_2rw
* cell instance $500 r0 *1 22.325,23.92
X$500 141 142 143 31 144 33 257 258 cell_2rw
* cell instance $501 r0 *1 23.5,23.92
X$501 145 146 147 31 148 33 257 258 cell_2rw
* cell instance $502 r0 *1 24.675,23.92
X$502 149 150 151 31 152 33 257 258 cell_2rw
* cell instance $503 r0 *1 25.85,23.92
X$503 153 154 155 31 156 33 257 258 cell_2rw
* cell instance $504 r0 *1 27.025,23.92
X$504 157 158 159 31 160 33 257 258 cell_2rw
* cell instance $505 r0 *1 28.2,23.92
X$505 161 162 163 31 164 33 257 258 cell_2rw
* cell instance $506 r0 *1 29.375,23.92
X$506 165 166 167 31 168 33 257 258 cell_2rw
* cell instance $507 r0 *1 30.55,23.92
X$507 169 170 171 31 172 33 257 258 cell_2rw
* cell instance $508 r0 *1 31.725,23.92
X$508 173 174 175 31 176 33 257 258 cell_2rw
* cell instance $509 r0 *1 32.9,23.92
X$509 177 178 179 31 180 33 257 258 cell_2rw
* cell instance $510 r0 *1 34.075,23.92
X$510 181 182 183 31 184 33 257 258 cell_2rw
* cell instance $511 r0 *1 35.25,23.92
X$511 185 186 187 31 188 33 257 258 cell_2rw
* cell instance $512 r0 *1 36.425,23.92
X$512 189 190 191 31 192 33 257 258 cell_2rw
* cell instance $513 m0 *1 1.175,26.91
X$513 65 66 67 34 68 32 257 258 cell_2rw
* cell instance $514 m0 *1 0,26.91
X$514 61 62 63 34 64 32 257 258 cell_2rw
* cell instance $515 m0 *1 2.35,26.91
X$515 69 70 71 34 72 32 257 258 cell_2rw
* cell instance $516 m0 *1 3.525,26.91
X$516 73 74 75 34 76 32 257 258 cell_2rw
* cell instance $517 m0 *1 4.7,26.91
X$517 77 78 79 34 80 32 257 258 cell_2rw
* cell instance $518 m0 *1 5.875,26.91
X$518 81 82 83 34 84 32 257 258 cell_2rw
* cell instance $519 m0 *1 7.05,26.91
X$519 85 86 87 34 88 32 257 258 cell_2rw
* cell instance $520 m0 *1 8.225,26.91
X$520 89 90 91 34 92 32 257 258 cell_2rw
* cell instance $521 m0 *1 9.4,26.91
X$521 93 94 95 34 96 32 257 258 cell_2rw
* cell instance $522 m0 *1 10.575,26.91
X$522 97 98 99 34 100 32 257 258 cell_2rw
* cell instance $523 m0 *1 11.75,26.91
X$523 101 102 103 34 104 32 257 258 cell_2rw
* cell instance $524 m0 *1 12.925,26.91
X$524 105 106 107 34 108 32 257 258 cell_2rw
* cell instance $525 m0 *1 14.1,26.91
X$525 109 110 111 34 112 32 257 258 cell_2rw
* cell instance $526 m0 *1 15.275,26.91
X$526 113 114 115 34 116 32 257 258 cell_2rw
* cell instance $527 m0 *1 16.45,26.91
X$527 117 118 119 34 120 32 257 258 cell_2rw
* cell instance $528 m0 *1 17.625,26.91
X$528 121 122 123 34 124 32 257 258 cell_2rw
* cell instance $529 m0 *1 18.8,26.91
X$529 129 130 131 34 132 32 257 258 cell_2rw
* cell instance $530 m0 *1 19.975,26.91
X$530 133 134 135 34 136 32 257 258 cell_2rw
* cell instance $531 m0 *1 21.15,26.91
X$531 137 138 139 34 140 32 257 258 cell_2rw
* cell instance $532 m0 *1 22.325,26.91
X$532 141 142 143 34 144 32 257 258 cell_2rw
* cell instance $533 m0 *1 23.5,26.91
X$533 145 146 147 34 148 32 257 258 cell_2rw
* cell instance $534 m0 *1 24.675,26.91
X$534 149 150 151 34 152 32 257 258 cell_2rw
* cell instance $535 m0 *1 25.85,26.91
X$535 153 154 155 34 156 32 257 258 cell_2rw
* cell instance $536 m0 *1 27.025,26.91
X$536 157 158 159 34 160 32 257 258 cell_2rw
* cell instance $537 m0 *1 28.2,26.91
X$537 161 162 163 34 164 32 257 258 cell_2rw
* cell instance $538 m0 *1 29.375,26.91
X$538 165 166 167 34 168 32 257 258 cell_2rw
* cell instance $539 m0 *1 30.55,26.91
X$539 169 170 171 34 172 32 257 258 cell_2rw
* cell instance $540 m0 *1 31.725,26.91
X$540 173 174 175 34 176 32 257 258 cell_2rw
* cell instance $541 m0 *1 32.9,26.91
X$541 177 178 179 34 180 32 257 258 cell_2rw
* cell instance $542 m0 *1 34.075,26.91
X$542 181 182 183 34 184 32 257 258 cell_2rw
* cell instance $543 m0 *1 35.25,26.91
X$543 185 186 187 34 188 32 257 258 cell_2rw
* cell instance $544 m0 *1 36.425,26.91
X$544 189 190 191 34 192 32 257 258 cell_2rw
* cell instance $545 m0 *1 1.175,23.92
X$545 65 66 67 35 68 36 257 258 cell_2rw
* cell instance $546 m0 *1 0,23.92
X$546 61 62 63 35 64 36 257 258 cell_2rw
* cell instance $547 m0 *1 2.35,23.92
X$547 69 70 71 35 72 36 257 258 cell_2rw
* cell instance $548 m0 *1 3.525,23.92
X$548 73 74 75 35 76 36 257 258 cell_2rw
* cell instance $549 m0 *1 4.7,23.92
X$549 77 78 79 35 80 36 257 258 cell_2rw
* cell instance $550 m0 *1 5.875,23.92
X$550 81 82 83 35 84 36 257 258 cell_2rw
* cell instance $551 m0 *1 7.05,23.92
X$551 85 86 87 35 88 36 257 258 cell_2rw
* cell instance $552 m0 *1 8.225,23.92
X$552 89 90 91 35 92 36 257 258 cell_2rw
* cell instance $553 m0 *1 9.4,23.92
X$553 93 94 95 35 96 36 257 258 cell_2rw
* cell instance $554 m0 *1 10.575,23.92
X$554 97 98 99 35 100 36 257 258 cell_2rw
* cell instance $555 m0 *1 11.75,23.92
X$555 101 102 103 35 104 36 257 258 cell_2rw
* cell instance $556 m0 *1 12.925,23.92
X$556 105 106 107 35 108 36 257 258 cell_2rw
* cell instance $557 m0 *1 14.1,23.92
X$557 109 110 111 35 112 36 257 258 cell_2rw
* cell instance $558 m0 *1 15.275,23.92
X$558 113 114 115 35 116 36 257 258 cell_2rw
* cell instance $559 m0 *1 16.45,23.92
X$559 117 118 119 35 120 36 257 258 cell_2rw
* cell instance $560 m0 *1 17.625,23.92
X$560 121 122 123 35 124 36 257 258 cell_2rw
* cell instance $561 m0 *1 18.8,23.92
X$561 129 130 131 35 132 36 257 258 cell_2rw
* cell instance $562 m0 *1 19.975,23.92
X$562 133 134 135 35 136 36 257 258 cell_2rw
* cell instance $563 m0 *1 21.15,23.92
X$563 137 138 139 35 140 36 257 258 cell_2rw
* cell instance $564 m0 *1 22.325,23.92
X$564 141 142 143 35 144 36 257 258 cell_2rw
* cell instance $565 m0 *1 23.5,23.92
X$565 145 146 147 35 148 36 257 258 cell_2rw
* cell instance $566 m0 *1 24.675,23.92
X$566 149 150 151 35 152 36 257 258 cell_2rw
* cell instance $567 m0 *1 25.85,23.92
X$567 153 154 155 35 156 36 257 258 cell_2rw
* cell instance $568 m0 *1 27.025,23.92
X$568 157 158 159 35 160 36 257 258 cell_2rw
* cell instance $569 m0 *1 28.2,23.92
X$569 161 162 163 35 164 36 257 258 cell_2rw
* cell instance $570 m0 *1 29.375,23.92
X$570 165 166 167 35 168 36 257 258 cell_2rw
* cell instance $571 m0 *1 30.55,23.92
X$571 169 170 171 35 172 36 257 258 cell_2rw
* cell instance $572 m0 *1 31.725,23.92
X$572 173 174 175 35 176 36 257 258 cell_2rw
* cell instance $573 m0 *1 32.9,23.92
X$573 177 178 179 35 180 36 257 258 cell_2rw
* cell instance $574 m0 *1 34.075,23.92
X$574 181 182 183 35 184 36 257 258 cell_2rw
* cell instance $575 m0 *1 35.25,23.92
X$575 185 186 187 35 188 36 257 258 cell_2rw
* cell instance $576 m0 *1 36.425,23.92
X$576 189 190 191 35 192 36 257 258 cell_2rw
* cell instance $577 r0 *1 1.175,29.9
X$577 65 66 67 37 68 38 257 258 cell_2rw
* cell instance $578 r0 *1 0,29.9
X$578 61 62 63 37 64 38 257 258 cell_2rw
* cell instance $579 r0 *1 2.35,29.9
X$579 69 70 71 37 72 38 257 258 cell_2rw
* cell instance $580 r0 *1 3.525,29.9
X$580 73 74 75 37 76 38 257 258 cell_2rw
* cell instance $581 r0 *1 4.7,29.9
X$581 77 78 79 37 80 38 257 258 cell_2rw
* cell instance $582 r0 *1 5.875,29.9
X$582 81 82 83 37 84 38 257 258 cell_2rw
* cell instance $583 r0 *1 7.05,29.9
X$583 85 86 87 37 88 38 257 258 cell_2rw
* cell instance $584 r0 *1 8.225,29.9
X$584 89 90 91 37 92 38 257 258 cell_2rw
* cell instance $585 r0 *1 9.4,29.9
X$585 93 94 95 37 96 38 257 258 cell_2rw
* cell instance $586 r0 *1 10.575,29.9
X$586 97 98 99 37 100 38 257 258 cell_2rw
* cell instance $587 r0 *1 11.75,29.9
X$587 101 102 103 37 104 38 257 258 cell_2rw
* cell instance $588 r0 *1 12.925,29.9
X$588 105 106 107 37 108 38 257 258 cell_2rw
* cell instance $589 r0 *1 14.1,29.9
X$589 109 110 111 37 112 38 257 258 cell_2rw
* cell instance $590 r0 *1 15.275,29.9
X$590 113 114 115 37 116 38 257 258 cell_2rw
* cell instance $591 r0 *1 16.45,29.9
X$591 117 118 119 37 120 38 257 258 cell_2rw
* cell instance $592 r0 *1 17.625,29.9
X$592 121 122 123 37 124 38 257 258 cell_2rw
* cell instance $593 r0 *1 18.8,29.9
X$593 129 130 131 37 132 38 257 258 cell_2rw
* cell instance $594 r0 *1 19.975,29.9
X$594 133 134 135 37 136 38 257 258 cell_2rw
* cell instance $595 r0 *1 21.15,29.9
X$595 137 138 139 37 140 38 257 258 cell_2rw
* cell instance $596 r0 *1 22.325,29.9
X$596 141 142 143 37 144 38 257 258 cell_2rw
* cell instance $597 r0 *1 23.5,29.9
X$597 145 146 147 37 148 38 257 258 cell_2rw
* cell instance $598 r0 *1 24.675,29.9
X$598 149 150 151 37 152 38 257 258 cell_2rw
* cell instance $599 r0 *1 25.85,29.9
X$599 153 154 155 37 156 38 257 258 cell_2rw
* cell instance $600 r0 *1 27.025,29.9
X$600 157 158 159 37 160 38 257 258 cell_2rw
* cell instance $601 r0 *1 28.2,29.9
X$601 161 162 163 37 164 38 257 258 cell_2rw
* cell instance $602 r0 *1 29.375,29.9
X$602 165 166 167 37 168 38 257 258 cell_2rw
* cell instance $603 r0 *1 30.55,29.9
X$603 169 170 171 37 172 38 257 258 cell_2rw
* cell instance $604 r0 *1 31.725,29.9
X$604 173 174 175 37 176 38 257 258 cell_2rw
* cell instance $605 r0 *1 32.9,29.9
X$605 177 178 179 37 180 38 257 258 cell_2rw
* cell instance $606 r0 *1 34.075,29.9
X$606 181 182 183 37 184 38 257 258 cell_2rw
* cell instance $607 r0 *1 35.25,29.9
X$607 185 186 187 37 188 38 257 258 cell_2rw
* cell instance $608 r0 *1 36.425,29.9
X$608 189 190 191 37 192 38 257 258 cell_2rw
* cell instance $609 r0 *1 1.175,26.91
X$609 65 66 67 42 68 39 257 258 cell_2rw
* cell instance $610 r0 *1 0,26.91
X$610 61 62 63 42 64 39 257 258 cell_2rw
* cell instance $611 r0 *1 2.35,26.91
X$611 69 70 71 42 72 39 257 258 cell_2rw
* cell instance $612 r0 *1 3.525,26.91
X$612 73 74 75 42 76 39 257 258 cell_2rw
* cell instance $613 r0 *1 4.7,26.91
X$613 77 78 79 42 80 39 257 258 cell_2rw
* cell instance $614 r0 *1 5.875,26.91
X$614 81 82 83 42 84 39 257 258 cell_2rw
* cell instance $615 r0 *1 7.05,26.91
X$615 85 86 87 42 88 39 257 258 cell_2rw
* cell instance $616 r0 *1 8.225,26.91
X$616 89 90 91 42 92 39 257 258 cell_2rw
* cell instance $617 r0 *1 9.4,26.91
X$617 93 94 95 42 96 39 257 258 cell_2rw
* cell instance $618 r0 *1 10.575,26.91
X$618 97 98 99 42 100 39 257 258 cell_2rw
* cell instance $619 r0 *1 11.75,26.91
X$619 101 102 103 42 104 39 257 258 cell_2rw
* cell instance $620 r0 *1 12.925,26.91
X$620 105 106 107 42 108 39 257 258 cell_2rw
* cell instance $621 r0 *1 14.1,26.91
X$621 109 110 111 42 112 39 257 258 cell_2rw
* cell instance $622 r0 *1 15.275,26.91
X$622 113 114 115 42 116 39 257 258 cell_2rw
* cell instance $623 r0 *1 16.45,26.91
X$623 117 118 119 42 120 39 257 258 cell_2rw
* cell instance $624 r0 *1 17.625,26.91
X$624 121 122 123 42 124 39 257 258 cell_2rw
* cell instance $625 r0 *1 18.8,26.91
X$625 129 130 131 42 132 39 257 258 cell_2rw
* cell instance $626 r0 *1 19.975,26.91
X$626 133 134 135 42 136 39 257 258 cell_2rw
* cell instance $627 r0 *1 21.15,26.91
X$627 137 138 139 42 140 39 257 258 cell_2rw
* cell instance $628 r0 *1 22.325,26.91
X$628 141 142 143 42 144 39 257 258 cell_2rw
* cell instance $629 r0 *1 23.5,26.91
X$629 145 146 147 42 148 39 257 258 cell_2rw
* cell instance $630 r0 *1 24.675,26.91
X$630 149 150 151 42 152 39 257 258 cell_2rw
* cell instance $631 r0 *1 25.85,26.91
X$631 153 154 155 42 156 39 257 258 cell_2rw
* cell instance $632 r0 *1 27.025,26.91
X$632 157 158 159 42 160 39 257 258 cell_2rw
* cell instance $633 r0 *1 28.2,26.91
X$633 161 162 163 42 164 39 257 258 cell_2rw
* cell instance $634 r0 *1 29.375,26.91
X$634 165 166 167 42 168 39 257 258 cell_2rw
* cell instance $635 r0 *1 30.55,26.91
X$635 169 170 171 42 172 39 257 258 cell_2rw
* cell instance $636 r0 *1 31.725,26.91
X$636 173 174 175 42 176 39 257 258 cell_2rw
* cell instance $637 r0 *1 32.9,26.91
X$637 177 178 179 42 180 39 257 258 cell_2rw
* cell instance $638 r0 *1 34.075,26.91
X$638 181 182 183 42 184 39 257 258 cell_2rw
* cell instance $639 r0 *1 35.25,26.91
X$639 185 186 187 42 188 39 257 258 cell_2rw
* cell instance $640 r0 *1 36.425,26.91
X$640 189 190 191 42 192 39 257 258 cell_2rw
* cell instance $641 m0 *1 1.175,29.9
X$641 65 66 67 41 68 40 257 258 cell_2rw
* cell instance $642 m0 *1 0,29.9
X$642 61 62 63 41 64 40 257 258 cell_2rw
* cell instance $643 m0 *1 2.35,29.9
X$643 69 70 71 41 72 40 257 258 cell_2rw
* cell instance $644 m0 *1 3.525,29.9
X$644 73 74 75 41 76 40 257 258 cell_2rw
* cell instance $645 m0 *1 4.7,29.9
X$645 77 78 79 41 80 40 257 258 cell_2rw
* cell instance $646 m0 *1 5.875,29.9
X$646 81 82 83 41 84 40 257 258 cell_2rw
* cell instance $647 m0 *1 7.05,29.9
X$647 85 86 87 41 88 40 257 258 cell_2rw
* cell instance $648 m0 *1 8.225,29.9
X$648 89 90 91 41 92 40 257 258 cell_2rw
* cell instance $649 m0 *1 9.4,29.9
X$649 93 94 95 41 96 40 257 258 cell_2rw
* cell instance $650 m0 *1 10.575,29.9
X$650 97 98 99 41 100 40 257 258 cell_2rw
* cell instance $651 m0 *1 11.75,29.9
X$651 101 102 103 41 104 40 257 258 cell_2rw
* cell instance $652 m0 *1 12.925,29.9
X$652 105 106 107 41 108 40 257 258 cell_2rw
* cell instance $653 m0 *1 14.1,29.9
X$653 109 110 111 41 112 40 257 258 cell_2rw
* cell instance $654 m0 *1 15.275,29.9
X$654 113 114 115 41 116 40 257 258 cell_2rw
* cell instance $655 m0 *1 16.45,29.9
X$655 117 118 119 41 120 40 257 258 cell_2rw
* cell instance $656 m0 *1 17.625,29.9
X$656 121 122 123 41 124 40 257 258 cell_2rw
* cell instance $657 m0 *1 18.8,29.9
X$657 129 130 131 41 132 40 257 258 cell_2rw
* cell instance $658 m0 *1 19.975,29.9
X$658 133 134 135 41 136 40 257 258 cell_2rw
* cell instance $659 m0 *1 21.15,29.9
X$659 137 138 139 41 140 40 257 258 cell_2rw
* cell instance $660 m0 *1 22.325,29.9
X$660 141 142 143 41 144 40 257 258 cell_2rw
* cell instance $661 m0 *1 23.5,29.9
X$661 145 146 147 41 148 40 257 258 cell_2rw
* cell instance $662 m0 *1 24.675,29.9
X$662 149 150 151 41 152 40 257 258 cell_2rw
* cell instance $663 m0 *1 25.85,29.9
X$663 153 154 155 41 156 40 257 258 cell_2rw
* cell instance $664 m0 *1 27.025,29.9
X$664 157 158 159 41 160 40 257 258 cell_2rw
* cell instance $665 m0 *1 28.2,29.9
X$665 161 162 163 41 164 40 257 258 cell_2rw
* cell instance $666 m0 *1 29.375,29.9
X$666 165 166 167 41 168 40 257 258 cell_2rw
* cell instance $667 m0 *1 30.55,29.9
X$667 169 170 171 41 172 40 257 258 cell_2rw
* cell instance $668 m0 *1 31.725,29.9
X$668 173 174 175 41 176 40 257 258 cell_2rw
* cell instance $669 m0 *1 32.9,29.9
X$669 177 178 179 41 180 40 257 258 cell_2rw
* cell instance $670 m0 *1 34.075,29.9
X$670 181 182 183 41 184 40 257 258 cell_2rw
* cell instance $671 m0 *1 35.25,29.9
X$671 185 186 187 41 188 40 257 258 cell_2rw
* cell instance $672 m0 *1 36.425,29.9
X$672 189 190 191 41 192 40 257 258 cell_2rw
* cell instance $673 r0 *1 1.175,32.89
X$673 65 66 67 44 68 43 257 258 cell_2rw
* cell instance $674 r0 *1 0,32.89
X$674 61 62 63 44 64 43 257 258 cell_2rw
* cell instance $675 r0 *1 2.35,32.89
X$675 69 70 71 44 72 43 257 258 cell_2rw
* cell instance $676 r0 *1 3.525,32.89
X$676 73 74 75 44 76 43 257 258 cell_2rw
* cell instance $677 r0 *1 4.7,32.89
X$677 77 78 79 44 80 43 257 258 cell_2rw
* cell instance $678 r0 *1 5.875,32.89
X$678 81 82 83 44 84 43 257 258 cell_2rw
* cell instance $679 r0 *1 7.05,32.89
X$679 85 86 87 44 88 43 257 258 cell_2rw
* cell instance $680 r0 *1 8.225,32.89
X$680 89 90 91 44 92 43 257 258 cell_2rw
* cell instance $681 r0 *1 9.4,32.89
X$681 93 94 95 44 96 43 257 258 cell_2rw
* cell instance $682 r0 *1 10.575,32.89
X$682 97 98 99 44 100 43 257 258 cell_2rw
* cell instance $683 r0 *1 11.75,32.89
X$683 101 102 103 44 104 43 257 258 cell_2rw
* cell instance $684 r0 *1 12.925,32.89
X$684 105 106 107 44 108 43 257 258 cell_2rw
* cell instance $685 r0 *1 14.1,32.89
X$685 109 110 111 44 112 43 257 258 cell_2rw
* cell instance $686 r0 *1 15.275,32.89
X$686 113 114 115 44 116 43 257 258 cell_2rw
* cell instance $687 r0 *1 16.45,32.89
X$687 117 118 119 44 120 43 257 258 cell_2rw
* cell instance $688 r0 *1 17.625,32.89
X$688 121 122 123 44 124 43 257 258 cell_2rw
* cell instance $689 r0 *1 18.8,32.89
X$689 129 130 131 44 132 43 257 258 cell_2rw
* cell instance $690 r0 *1 19.975,32.89
X$690 133 134 135 44 136 43 257 258 cell_2rw
* cell instance $691 r0 *1 21.15,32.89
X$691 137 138 139 44 140 43 257 258 cell_2rw
* cell instance $692 r0 *1 22.325,32.89
X$692 141 142 143 44 144 43 257 258 cell_2rw
* cell instance $693 r0 *1 23.5,32.89
X$693 145 146 147 44 148 43 257 258 cell_2rw
* cell instance $694 r0 *1 24.675,32.89
X$694 149 150 151 44 152 43 257 258 cell_2rw
* cell instance $695 r0 *1 25.85,32.89
X$695 153 154 155 44 156 43 257 258 cell_2rw
* cell instance $696 r0 *1 27.025,32.89
X$696 157 158 159 44 160 43 257 258 cell_2rw
* cell instance $697 r0 *1 28.2,32.89
X$697 161 162 163 44 164 43 257 258 cell_2rw
* cell instance $698 r0 *1 29.375,32.89
X$698 165 166 167 44 168 43 257 258 cell_2rw
* cell instance $699 r0 *1 30.55,32.89
X$699 169 170 171 44 172 43 257 258 cell_2rw
* cell instance $700 r0 *1 31.725,32.89
X$700 173 174 175 44 176 43 257 258 cell_2rw
* cell instance $701 r0 *1 32.9,32.89
X$701 177 178 179 44 180 43 257 258 cell_2rw
* cell instance $702 r0 *1 34.075,32.89
X$702 181 182 183 44 184 43 257 258 cell_2rw
* cell instance $703 r0 *1 35.25,32.89
X$703 185 186 187 44 188 43 257 258 cell_2rw
* cell instance $704 r0 *1 36.425,32.89
X$704 189 190 191 44 192 43 257 258 cell_2rw
* cell instance $705 m0 *1 1.175,35.88
X$705 65 66 67 45 68 46 257 258 cell_2rw
* cell instance $706 m0 *1 0,35.88
X$706 61 62 63 45 64 46 257 258 cell_2rw
* cell instance $707 m0 *1 2.35,35.88
X$707 69 70 71 45 72 46 257 258 cell_2rw
* cell instance $708 m0 *1 3.525,35.88
X$708 73 74 75 45 76 46 257 258 cell_2rw
* cell instance $709 m0 *1 4.7,35.88
X$709 77 78 79 45 80 46 257 258 cell_2rw
* cell instance $710 m0 *1 5.875,35.88
X$710 81 82 83 45 84 46 257 258 cell_2rw
* cell instance $711 m0 *1 7.05,35.88
X$711 85 86 87 45 88 46 257 258 cell_2rw
* cell instance $712 m0 *1 8.225,35.88
X$712 89 90 91 45 92 46 257 258 cell_2rw
* cell instance $713 m0 *1 9.4,35.88
X$713 93 94 95 45 96 46 257 258 cell_2rw
* cell instance $714 m0 *1 10.575,35.88
X$714 97 98 99 45 100 46 257 258 cell_2rw
* cell instance $715 m0 *1 11.75,35.88
X$715 101 102 103 45 104 46 257 258 cell_2rw
* cell instance $716 m0 *1 12.925,35.88
X$716 105 106 107 45 108 46 257 258 cell_2rw
* cell instance $717 m0 *1 14.1,35.88
X$717 109 110 111 45 112 46 257 258 cell_2rw
* cell instance $718 m0 *1 15.275,35.88
X$718 113 114 115 45 116 46 257 258 cell_2rw
* cell instance $719 m0 *1 16.45,35.88
X$719 117 118 119 45 120 46 257 258 cell_2rw
* cell instance $720 m0 *1 17.625,35.88
X$720 121 122 123 45 124 46 257 258 cell_2rw
* cell instance $721 m0 *1 18.8,35.88
X$721 129 130 131 45 132 46 257 258 cell_2rw
* cell instance $722 m0 *1 19.975,35.88
X$722 133 134 135 45 136 46 257 258 cell_2rw
* cell instance $723 m0 *1 21.15,35.88
X$723 137 138 139 45 140 46 257 258 cell_2rw
* cell instance $724 m0 *1 22.325,35.88
X$724 141 142 143 45 144 46 257 258 cell_2rw
* cell instance $725 m0 *1 23.5,35.88
X$725 145 146 147 45 148 46 257 258 cell_2rw
* cell instance $726 m0 *1 24.675,35.88
X$726 149 150 151 45 152 46 257 258 cell_2rw
* cell instance $727 m0 *1 25.85,35.88
X$727 153 154 155 45 156 46 257 258 cell_2rw
* cell instance $728 m0 *1 27.025,35.88
X$728 157 158 159 45 160 46 257 258 cell_2rw
* cell instance $729 m0 *1 28.2,35.88
X$729 161 162 163 45 164 46 257 258 cell_2rw
* cell instance $730 m0 *1 29.375,35.88
X$730 165 166 167 45 168 46 257 258 cell_2rw
* cell instance $731 m0 *1 30.55,35.88
X$731 169 170 171 45 172 46 257 258 cell_2rw
* cell instance $732 m0 *1 31.725,35.88
X$732 173 174 175 45 176 46 257 258 cell_2rw
* cell instance $733 m0 *1 32.9,35.88
X$733 177 178 179 45 180 46 257 258 cell_2rw
* cell instance $734 m0 *1 34.075,35.88
X$734 181 182 183 45 184 46 257 258 cell_2rw
* cell instance $735 m0 *1 35.25,35.88
X$735 185 186 187 45 188 46 257 258 cell_2rw
* cell instance $736 m0 *1 36.425,35.88
X$736 189 190 191 45 192 46 257 258 cell_2rw
* cell instance $737 m0 *1 1.175,32.89
X$737 65 66 67 48 68 47 257 258 cell_2rw
* cell instance $738 m0 *1 0,32.89
X$738 61 62 63 48 64 47 257 258 cell_2rw
* cell instance $739 m0 *1 2.35,32.89
X$739 69 70 71 48 72 47 257 258 cell_2rw
* cell instance $740 m0 *1 3.525,32.89
X$740 73 74 75 48 76 47 257 258 cell_2rw
* cell instance $741 m0 *1 4.7,32.89
X$741 77 78 79 48 80 47 257 258 cell_2rw
* cell instance $742 m0 *1 5.875,32.89
X$742 81 82 83 48 84 47 257 258 cell_2rw
* cell instance $743 m0 *1 7.05,32.89
X$743 85 86 87 48 88 47 257 258 cell_2rw
* cell instance $744 m0 *1 8.225,32.89
X$744 89 90 91 48 92 47 257 258 cell_2rw
* cell instance $745 m0 *1 9.4,32.89
X$745 93 94 95 48 96 47 257 258 cell_2rw
* cell instance $746 m0 *1 10.575,32.89
X$746 97 98 99 48 100 47 257 258 cell_2rw
* cell instance $747 m0 *1 11.75,32.89
X$747 101 102 103 48 104 47 257 258 cell_2rw
* cell instance $748 m0 *1 12.925,32.89
X$748 105 106 107 48 108 47 257 258 cell_2rw
* cell instance $749 m0 *1 14.1,32.89
X$749 109 110 111 48 112 47 257 258 cell_2rw
* cell instance $750 m0 *1 15.275,32.89
X$750 113 114 115 48 116 47 257 258 cell_2rw
* cell instance $751 m0 *1 16.45,32.89
X$751 117 118 119 48 120 47 257 258 cell_2rw
* cell instance $752 m0 *1 17.625,32.89
X$752 121 122 123 48 124 47 257 258 cell_2rw
* cell instance $753 m0 *1 18.8,32.89
X$753 129 130 131 48 132 47 257 258 cell_2rw
* cell instance $754 m0 *1 19.975,32.89
X$754 133 134 135 48 136 47 257 258 cell_2rw
* cell instance $755 m0 *1 21.15,32.89
X$755 137 138 139 48 140 47 257 258 cell_2rw
* cell instance $756 m0 *1 22.325,32.89
X$756 141 142 143 48 144 47 257 258 cell_2rw
* cell instance $757 m0 *1 23.5,32.89
X$757 145 146 147 48 148 47 257 258 cell_2rw
* cell instance $758 m0 *1 24.675,32.89
X$758 149 150 151 48 152 47 257 258 cell_2rw
* cell instance $759 m0 *1 25.85,32.89
X$759 153 154 155 48 156 47 257 258 cell_2rw
* cell instance $760 m0 *1 27.025,32.89
X$760 157 158 159 48 160 47 257 258 cell_2rw
* cell instance $761 m0 *1 28.2,32.89
X$761 161 162 163 48 164 47 257 258 cell_2rw
* cell instance $762 m0 *1 29.375,32.89
X$762 165 166 167 48 168 47 257 258 cell_2rw
* cell instance $763 m0 *1 30.55,32.89
X$763 169 170 171 48 172 47 257 258 cell_2rw
* cell instance $764 m0 *1 31.725,32.89
X$764 173 174 175 48 176 47 257 258 cell_2rw
* cell instance $765 m0 *1 32.9,32.89
X$765 177 178 179 48 180 47 257 258 cell_2rw
* cell instance $766 m0 *1 34.075,32.89
X$766 181 182 183 48 184 47 257 258 cell_2rw
* cell instance $767 m0 *1 35.25,32.89
X$767 185 186 187 48 188 47 257 258 cell_2rw
* cell instance $768 m0 *1 36.425,32.89
X$768 189 190 191 48 192 47 257 258 cell_2rw
* cell instance $769 m0 *1 1.175,38.87
X$769 65 66 67 54 68 49 257 258 cell_2rw
* cell instance $770 m0 *1 0,38.87
X$770 61 62 63 54 64 49 257 258 cell_2rw
* cell instance $771 m0 *1 2.35,38.87
X$771 69 70 71 54 72 49 257 258 cell_2rw
* cell instance $772 m0 *1 3.525,38.87
X$772 73 74 75 54 76 49 257 258 cell_2rw
* cell instance $773 m0 *1 4.7,38.87
X$773 77 78 79 54 80 49 257 258 cell_2rw
* cell instance $774 m0 *1 5.875,38.87
X$774 81 82 83 54 84 49 257 258 cell_2rw
* cell instance $775 m0 *1 7.05,38.87
X$775 85 86 87 54 88 49 257 258 cell_2rw
* cell instance $776 m0 *1 8.225,38.87
X$776 89 90 91 54 92 49 257 258 cell_2rw
* cell instance $777 m0 *1 9.4,38.87
X$777 93 94 95 54 96 49 257 258 cell_2rw
* cell instance $778 m0 *1 10.575,38.87
X$778 97 98 99 54 100 49 257 258 cell_2rw
* cell instance $779 m0 *1 11.75,38.87
X$779 101 102 103 54 104 49 257 258 cell_2rw
* cell instance $780 m0 *1 12.925,38.87
X$780 105 106 107 54 108 49 257 258 cell_2rw
* cell instance $781 m0 *1 14.1,38.87
X$781 109 110 111 54 112 49 257 258 cell_2rw
* cell instance $782 m0 *1 15.275,38.87
X$782 113 114 115 54 116 49 257 258 cell_2rw
* cell instance $783 m0 *1 16.45,38.87
X$783 117 118 119 54 120 49 257 258 cell_2rw
* cell instance $784 m0 *1 17.625,38.87
X$784 121 122 123 54 124 49 257 258 cell_2rw
* cell instance $785 m0 *1 18.8,38.87
X$785 129 130 131 54 132 49 257 258 cell_2rw
* cell instance $786 m0 *1 19.975,38.87
X$786 133 134 135 54 136 49 257 258 cell_2rw
* cell instance $787 m0 *1 21.15,38.87
X$787 137 138 139 54 140 49 257 258 cell_2rw
* cell instance $788 m0 *1 22.325,38.87
X$788 141 142 143 54 144 49 257 258 cell_2rw
* cell instance $789 m0 *1 23.5,38.87
X$789 145 146 147 54 148 49 257 258 cell_2rw
* cell instance $790 m0 *1 24.675,38.87
X$790 149 150 151 54 152 49 257 258 cell_2rw
* cell instance $791 m0 *1 25.85,38.87
X$791 153 154 155 54 156 49 257 258 cell_2rw
* cell instance $792 m0 *1 27.025,38.87
X$792 157 158 159 54 160 49 257 258 cell_2rw
* cell instance $793 m0 *1 28.2,38.87
X$793 161 162 163 54 164 49 257 258 cell_2rw
* cell instance $794 m0 *1 29.375,38.87
X$794 165 166 167 54 168 49 257 258 cell_2rw
* cell instance $795 m0 *1 30.55,38.87
X$795 169 170 171 54 172 49 257 258 cell_2rw
* cell instance $796 m0 *1 31.725,38.87
X$796 173 174 175 54 176 49 257 258 cell_2rw
* cell instance $797 m0 *1 32.9,38.87
X$797 177 178 179 54 180 49 257 258 cell_2rw
* cell instance $798 m0 *1 34.075,38.87
X$798 181 182 183 54 184 49 257 258 cell_2rw
* cell instance $799 m0 *1 35.25,38.87
X$799 185 186 187 54 188 49 257 258 cell_2rw
* cell instance $800 m0 *1 36.425,38.87
X$800 189 190 191 54 192 49 257 258 cell_2rw
* cell instance $801 r0 *1 1.175,38.87
X$801 65 66 67 51 68 50 257 258 cell_2rw
* cell instance $802 r0 *1 0,38.87
X$802 61 62 63 51 64 50 257 258 cell_2rw
* cell instance $803 r0 *1 2.35,38.87
X$803 69 70 71 51 72 50 257 258 cell_2rw
* cell instance $804 r0 *1 3.525,38.87
X$804 73 74 75 51 76 50 257 258 cell_2rw
* cell instance $805 r0 *1 4.7,38.87
X$805 77 78 79 51 80 50 257 258 cell_2rw
* cell instance $806 r0 *1 5.875,38.87
X$806 81 82 83 51 84 50 257 258 cell_2rw
* cell instance $807 r0 *1 7.05,38.87
X$807 85 86 87 51 88 50 257 258 cell_2rw
* cell instance $808 r0 *1 8.225,38.87
X$808 89 90 91 51 92 50 257 258 cell_2rw
* cell instance $809 r0 *1 9.4,38.87
X$809 93 94 95 51 96 50 257 258 cell_2rw
* cell instance $810 r0 *1 10.575,38.87
X$810 97 98 99 51 100 50 257 258 cell_2rw
* cell instance $811 r0 *1 11.75,38.87
X$811 101 102 103 51 104 50 257 258 cell_2rw
* cell instance $812 r0 *1 12.925,38.87
X$812 105 106 107 51 108 50 257 258 cell_2rw
* cell instance $813 r0 *1 14.1,38.87
X$813 109 110 111 51 112 50 257 258 cell_2rw
* cell instance $814 r0 *1 15.275,38.87
X$814 113 114 115 51 116 50 257 258 cell_2rw
* cell instance $815 r0 *1 16.45,38.87
X$815 117 118 119 51 120 50 257 258 cell_2rw
* cell instance $816 r0 *1 17.625,38.87
X$816 121 122 123 51 124 50 257 258 cell_2rw
* cell instance $817 r0 *1 18.8,38.87
X$817 129 130 131 51 132 50 257 258 cell_2rw
* cell instance $818 r0 *1 19.975,38.87
X$818 133 134 135 51 136 50 257 258 cell_2rw
* cell instance $819 r0 *1 21.15,38.87
X$819 137 138 139 51 140 50 257 258 cell_2rw
* cell instance $820 r0 *1 22.325,38.87
X$820 141 142 143 51 144 50 257 258 cell_2rw
* cell instance $821 r0 *1 23.5,38.87
X$821 145 146 147 51 148 50 257 258 cell_2rw
* cell instance $822 r0 *1 24.675,38.87
X$822 149 150 151 51 152 50 257 258 cell_2rw
* cell instance $823 r0 *1 25.85,38.87
X$823 153 154 155 51 156 50 257 258 cell_2rw
* cell instance $824 r0 *1 27.025,38.87
X$824 157 158 159 51 160 50 257 258 cell_2rw
* cell instance $825 r0 *1 28.2,38.87
X$825 161 162 163 51 164 50 257 258 cell_2rw
* cell instance $826 r0 *1 29.375,38.87
X$826 165 166 167 51 168 50 257 258 cell_2rw
* cell instance $827 r0 *1 30.55,38.87
X$827 169 170 171 51 172 50 257 258 cell_2rw
* cell instance $828 r0 *1 31.725,38.87
X$828 173 174 175 51 176 50 257 258 cell_2rw
* cell instance $829 r0 *1 32.9,38.87
X$829 177 178 179 51 180 50 257 258 cell_2rw
* cell instance $830 r0 *1 34.075,38.87
X$830 181 182 183 51 184 50 257 258 cell_2rw
* cell instance $831 r0 *1 35.25,38.87
X$831 185 186 187 51 188 50 257 258 cell_2rw
* cell instance $832 r0 *1 36.425,38.87
X$832 189 190 191 51 192 50 257 258 cell_2rw
* cell instance $833 r0 *1 1.175,35.88
X$833 65 66 67 53 68 52 257 258 cell_2rw
* cell instance $834 r0 *1 0,35.88
X$834 61 62 63 53 64 52 257 258 cell_2rw
* cell instance $835 r0 *1 2.35,35.88
X$835 69 70 71 53 72 52 257 258 cell_2rw
* cell instance $836 r0 *1 3.525,35.88
X$836 73 74 75 53 76 52 257 258 cell_2rw
* cell instance $837 r0 *1 4.7,35.88
X$837 77 78 79 53 80 52 257 258 cell_2rw
* cell instance $838 r0 *1 5.875,35.88
X$838 81 82 83 53 84 52 257 258 cell_2rw
* cell instance $839 r0 *1 7.05,35.88
X$839 85 86 87 53 88 52 257 258 cell_2rw
* cell instance $840 r0 *1 8.225,35.88
X$840 89 90 91 53 92 52 257 258 cell_2rw
* cell instance $841 r0 *1 9.4,35.88
X$841 93 94 95 53 96 52 257 258 cell_2rw
* cell instance $842 r0 *1 10.575,35.88
X$842 97 98 99 53 100 52 257 258 cell_2rw
* cell instance $843 r0 *1 11.75,35.88
X$843 101 102 103 53 104 52 257 258 cell_2rw
* cell instance $844 r0 *1 12.925,35.88
X$844 105 106 107 53 108 52 257 258 cell_2rw
* cell instance $845 r0 *1 14.1,35.88
X$845 109 110 111 53 112 52 257 258 cell_2rw
* cell instance $846 r0 *1 15.275,35.88
X$846 113 114 115 53 116 52 257 258 cell_2rw
* cell instance $847 r0 *1 16.45,35.88
X$847 117 118 119 53 120 52 257 258 cell_2rw
* cell instance $848 r0 *1 17.625,35.88
X$848 121 122 123 53 124 52 257 258 cell_2rw
* cell instance $849 r0 *1 18.8,35.88
X$849 129 130 131 53 132 52 257 258 cell_2rw
* cell instance $850 r0 *1 19.975,35.88
X$850 133 134 135 53 136 52 257 258 cell_2rw
* cell instance $851 r0 *1 21.15,35.88
X$851 137 138 139 53 140 52 257 258 cell_2rw
* cell instance $852 r0 *1 22.325,35.88
X$852 141 142 143 53 144 52 257 258 cell_2rw
* cell instance $853 r0 *1 23.5,35.88
X$853 145 146 147 53 148 52 257 258 cell_2rw
* cell instance $854 r0 *1 24.675,35.88
X$854 149 150 151 53 152 52 257 258 cell_2rw
* cell instance $855 r0 *1 25.85,35.88
X$855 153 154 155 53 156 52 257 258 cell_2rw
* cell instance $856 r0 *1 27.025,35.88
X$856 157 158 159 53 160 52 257 258 cell_2rw
* cell instance $857 r0 *1 28.2,35.88
X$857 161 162 163 53 164 52 257 258 cell_2rw
* cell instance $858 r0 *1 29.375,35.88
X$858 165 166 167 53 168 52 257 258 cell_2rw
* cell instance $859 r0 *1 30.55,35.88
X$859 169 170 171 53 172 52 257 258 cell_2rw
* cell instance $860 r0 *1 31.725,35.88
X$860 173 174 175 53 176 52 257 258 cell_2rw
* cell instance $861 r0 *1 32.9,35.88
X$861 177 178 179 53 180 52 257 258 cell_2rw
* cell instance $862 r0 *1 34.075,35.88
X$862 181 182 183 53 184 52 257 258 cell_2rw
* cell instance $863 r0 *1 35.25,35.88
X$863 185 186 187 53 188 52 257 258 cell_2rw
* cell instance $864 r0 *1 36.425,35.88
X$864 189 190 191 53 192 52 257 258 cell_2rw
* cell instance $865 r0 *1 1.175,41.86
X$865 65 66 67 56 68 55 257 258 cell_2rw
* cell instance $866 r0 *1 0,41.86
X$866 61 62 63 56 64 55 257 258 cell_2rw
* cell instance $867 r0 *1 2.35,41.86
X$867 69 70 71 56 72 55 257 258 cell_2rw
* cell instance $868 r0 *1 3.525,41.86
X$868 73 74 75 56 76 55 257 258 cell_2rw
* cell instance $869 r0 *1 4.7,41.86
X$869 77 78 79 56 80 55 257 258 cell_2rw
* cell instance $870 r0 *1 5.875,41.86
X$870 81 82 83 56 84 55 257 258 cell_2rw
* cell instance $871 r0 *1 7.05,41.86
X$871 85 86 87 56 88 55 257 258 cell_2rw
* cell instance $872 r0 *1 8.225,41.86
X$872 89 90 91 56 92 55 257 258 cell_2rw
* cell instance $873 r0 *1 9.4,41.86
X$873 93 94 95 56 96 55 257 258 cell_2rw
* cell instance $874 r0 *1 10.575,41.86
X$874 97 98 99 56 100 55 257 258 cell_2rw
* cell instance $875 r0 *1 11.75,41.86
X$875 101 102 103 56 104 55 257 258 cell_2rw
* cell instance $876 r0 *1 12.925,41.86
X$876 105 106 107 56 108 55 257 258 cell_2rw
* cell instance $877 r0 *1 14.1,41.86
X$877 109 110 111 56 112 55 257 258 cell_2rw
* cell instance $878 r0 *1 15.275,41.86
X$878 113 114 115 56 116 55 257 258 cell_2rw
* cell instance $879 r0 *1 16.45,41.86
X$879 117 118 119 56 120 55 257 258 cell_2rw
* cell instance $880 r0 *1 17.625,41.86
X$880 121 122 123 56 124 55 257 258 cell_2rw
* cell instance $881 r0 *1 18.8,41.86
X$881 129 130 131 56 132 55 257 258 cell_2rw
* cell instance $882 r0 *1 19.975,41.86
X$882 133 134 135 56 136 55 257 258 cell_2rw
* cell instance $883 r0 *1 21.15,41.86
X$883 137 138 139 56 140 55 257 258 cell_2rw
* cell instance $884 r0 *1 22.325,41.86
X$884 141 142 143 56 144 55 257 258 cell_2rw
* cell instance $885 r0 *1 23.5,41.86
X$885 145 146 147 56 148 55 257 258 cell_2rw
* cell instance $886 r0 *1 24.675,41.86
X$886 149 150 151 56 152 55 257 258 cell_2rw
* cell instance $887 r0 *1 25.85,41.86
X$887 153 154 155 56 156 55 257 258 cell_2rw
* cell instance $888 r0 *1 27.025,41.86
X$888 157 158 159 56 160 55 257 258 cell_2rw
* cell instance $889 r0 *1 28.2,41.86
X$889 161 162 163 56 164 55 257 258 cell_2rw
* cell instance $890 r0 *1 29.375,41.86
X$890 165 166 167 56 168 55 257 258 cell_2rw
* cell instance $891 r0 *1 30.55,41.86
X$891 169 170 171 56 172 55 257 258 cell_2rw
* cell instance $892 r0 *1 31.725,41.86
X$892 173 174 175 56 176 55 257 258 cell_2rw
* cell instance $893 r0 *1 32.9,41.86
X$893 177 178 179 56 180 55 257 258 cell_2rw
* cell instance $894 r0 *1 34.075,41.86
X$894 181 182 183 56 184 55 257 258 cell_2rw
* cell instance $895 r0 *1 35.25,41.86
X$895 185 186 187 56 188 55 257 258 cell_2rw
* cell instance $896 r0 *1 36.425,41.86
X$896 189 190 191 56 192 55 257 258 cell_2rw
* cell instance $897 m0 *1 1.175,44.85
X$897 65 66 67 60 68 57 257 258 cell_2rw
* cell instance $898 m0 *1 0,44.85
X$898 61 62 63 60 64 57 257 258 cell_2rw
* cell instance $899 m0 *1 2.35,44.85
X$899 69 70 71 60 72 57 257 258 cell_2rw
* cell instance $900 m0 *1 3.525,44.85
X$900 73 74 75 60 76 57 257 258 cell_2rw
* cell instance $901 m0 *1 4.7,44.85
X$901 77 78 79 60 80 57 257 258 cell_2rw
* cell instance $902 m0 *1 5.875,44.85
X$902 81 82 83 60 84 57 257 258 cell_2rw
* cell instance $903 m0 *1 7.05,44.85
X$903 85 86 87 60 88 57 257 258 cell_2rw
* cell instance $904 m0 *1 8.225,44.85
X$904 89 90 91 60 92 57 257 258 cell_2rw
* cell instance $905 m0 *1 9.4,44.85
X$905 93 94 95 60 96 57 257 258 cell_2rw
* cell instance $906 m0 *1 10.575,44.85
X$906 97 98 99 60 100 57 257 258 cell_2rw
* cell instance $907 m0 *1 11.75,44.85
X$907 101 102 103 60 104 57 257 258 cell_2rw
* cell instance $908 m0 *1 12.925,44.85
X$908 105 106 107 60 108 57 257 258 cell_2rw
* cell instance $909 m0 *1 14.1,44.85
X$909 109 110 111 60 112 57 257 258 cell_2rw
* cell instance $910 m0 *1 15.275,44.85
X$910 113 114 115 60 116 57 257 258 cell_2rw
* cell instance $911 m0 *1 16.45,44.85
X$911 117 118 119 60 120 57 257 258 cell_2rw
* cell instance $912 m0 *1 17.625,44.85
X$912 121 122 123 60 124 57 257 258 cell_2rw
* cell instance $913 m0 *1 18.8,44.85
X$913 129 130 131 60 132 57 257 258 cell_2rw
* cell instance $914 m0 *1 19.975,44.85
X$914 133 134 135 60 136 57 257 258 cell_2rw
* cell instance $915 m0 *1 21.15,44.85
X$915 137 138 139 60 140 57 257 258 cell_2rw
* cell instance $916 m0 *1 22.325,44.85
X$916 141 142 143 60 144 57 257 258 cell_2rw
* cell instance $917 m0 *1 23.5,44.85
X$917 145 146 147 60 148 57 257 258 cell_2rw
* cell instance $918 m0 *1 24.675,44.85
X$918 149 150 151 60 152 57 257 258 cell_2rw
* cell instance $919 m0 *1 25.85,44.85
X$919 153 154 155 60 156 57 257 258 cell_2rw
* cell instance $920 m0 *1 27.025,44.85
X$920 157 158 159 60 160 57 257 258 cell_2rw
* cell instance $921 m0 *1 28.2,44.85
X$921 161 162 163 60 164 57 257 258 cell_2rw
* cell instance $922 m0 *1 29.375,44.85
X$922 165 166 167 60 168 57 257 258 cell_2rw
* cell instance $923 m0 *1 30.55,44.85
X$923 169 170 171 60 172 57 257 258 cell_2rw
* cell instance $924 m0 *1 31.725,44.85
X$924 173 174 175 60 176 57 257 258 cell_2rw
* cell instance $925 m0 *1 32.9,44.85
X$925 177 178 179 60 180 57 257 258 cell_2rw
* cell instance $926 m0 *1 34.075,44.85
X$926 181 182 183 60 184 57 257 258 cell_2rw
* cell instance $927 m0 *1 35.25,44.85
X$927 185 186 187 60 188 57 257 258 cell_2rw
* cell instance $928 m0 *1 36.425,44.85
X$928 189 190 191 60 192 57 257 258 cell_2rw
* cell instance $929 m0 *1 1.175,41.86
X$929 65 66 67 59 68 58 257 258 cell_2rw
* cell instance $930 m0 *1 0,41.86
X$930 61 62 63 59 64 58 257 258 cell_2rw
* cell instance $931 m0 *1 2.35,41.86
X$931 69 70 71 59 72 58 257 258 cell_2rw
* cell instance $932 m0 *1 3.525,41.86
X$932 73 74 75 59 76 58 257 258 cell_2rw
* cell instance $933 m0 *1 4.7,41.86
X$933 77 78 79 59 80 58 257 258 cell_2rw
* cell instance $934 m0 *1 5.875,41.86
X$934 81 82 83 59 84 58 257 258 cell_2rw
* cell instance $935 m0 *1 7.05,41.86
X$935 85 86 87 59 88 58 257 258 cell_2rw
* cell instance $936 m0 *1 8.225,41.86
X$936 89 90 91 59 92 58 257 258 cell_2rw
* cell instance $937 m0 *1 9.4,41.86
X$937 93 94 95 59 96 58 257 258 cell_2rw
* cell instance $938 m0 *1 10.575,41.86
X$938 97 98 99 59 100 58 257 258 cell_2rw
* cell instance $939 m0 *1 11.75,41.86
X$939 101 102 103 59 104 58 257 258 cell_2rw
* cell instance $940 m0 *1 12.925,41.86
X$940 105 106 107 59 108 58 257 258 cell_2rw
* cell instance $941 m0 *1 14.1,41.86
X$941 109 110 111 59 112 58 257 258 cell_2rw
* cell instance $942 m0 *1 15.275,41.86
X$942 113 114 115 59 116 58 257 258 cell_2rw
* cell instance $943 m0 *1 16.45,41.86
X$943 117 118 119 59 120 58 257 258 cell_2rw
* cell instance $944 m0 *1 17.625,41.86
X$944 121 122 123 59 124 58 257 258 cell_2rw
* cell instance $945 m0 *1 18.8,41.86
X$945 129 130 131 59 132 58 257 258 cell_2rw
* cell instance $946 m0 *1 19.975,41.86
X$946 133 134 135 59 136 58 257 258 cell_2rw
* cell instance $947 m0 *1 21.15,41.86
X$947 137 138 139 59 140 58 257 258 cell_2rw
* cell instance $948 m0 *1 22.325,41.86
X$948 141 142 143 59 144 58 257 258 cell_2rw
* cell instance $949 m0 *1 23.5,41.86
X$949 145 146 147 59 148 58 257 258 cell_2rw
* cell instance $950 m0 *1 24.675,41.86
X$950 149 150 151 59 152 58 257 258 cell_2rw
* cell instance $951 m0 *1 25.85,41.86
X$951 153 154 155 59 156 58 257 258 cell_2rw
* cell instance $952 m0 *1 27.025,41.86
X$952 157 158 159 59 160 58 257 258 cell_2rw
* cell instance $953 m0 *1 28.2,41.86
X$953 161 162 163 59 164 58 257 258 cell_2rw
* cell instance $954 m0 *1 29.375,41.86
X$954 165 166 167 59 168 58 257 258 cell_2rw
* cell instance $955 m0 *1 30.55,41.86
X$955 169 170 171 59 172 58 257 258 cell_2rw
* cell instance $956 m0 *1 31.725,41.86
X$956 173 174 175 59 176 58 257 258 cell_2rw
* cell instance $957 m0 *1 32.9,41.86
X$957 177 178 179 59 180 58 257 258 cell_2rw
* cell instance $958 m0 *1 34.075,41.86
X$958 181 182 183 59 184 58 257 258 cell_2rw
* cell instance $959 m0 *1 35.25,41.86
X$959 185 186 187 59 188 58 257 258 cell_2rw
* cell instance $960 m0 *1 36.425,41.86
X$960 189 190 191 59 192 58 257 258 cell_2rw
* cell instance $961 r0 *1 0,44.85
X$961 61 62 63 127 64 128 257 258 cell_2rw
* cell instance $962 m0 *1 0,47.84
X$962 61 62 63 126 64 125 257 258 cell_2rw
* cell instance $963 m0 *1 0,50.83
X$963 61 62 63 195 64 197 257 258 cell_2rw
* cell instance $964 r0 *1 0,47.84
X$964 61 62 63 199 64 201 257 258 cell_2rw
* cell instance $965 r0 *1 0,50.83
X$965 61 62 63 202 64 194 257 258 cell_2rw
* cell instance $966 m0 *1 0,53.82
X$966 61 62 63 198 64 193 257 258 cell_2rw
* cell instance $967 r0 *1 0,53.82
X$967 61 62 63 196 64 200 257 258 cell_2rw
* cell instance $968 m0 *1 0,56.81
X$968 61 62 63 203 64 207 257 258 cell_2rw
* cell instance $969 r0 *1 0,56.81
X$969 61 62 63 206 64 208 257 258 cell_2rw
* cell instance $970 m0 *1 0,59.8
X$970 61 62 63 205 64 204 257 258 cell_2rw
* cell instance $971 r0 *1 0,59.8
X$971 61 62 63 214 64 213 257 258 cell_2rw
* cell instance $972 m0 *1 0,62.79
X$972 61 62 63 212 64 211 257 258 cell_2rw
* cell instance $973 r0 *1 0,62.79
X$973 61 62 63 210 64 209 257 258 cell_2rw
* cell instance $974 m0 *1 0,65.78
X$974 61 62 63 219 64 217 257 258 cell_2rw
* cell instance $975 r0 *1 0,65.78
X$975 61 62 63 216 64 215 257 258 cell_2rw
* cell instance $976 m0 *1 0,68.77
X$976 61 62 63 218 64 220 257 258 cell_2rw
* cell instance $977 r0 *1 0,68.77
X$977 61 62 63 224 64 223 257 258 cell_2rw
* cell instance $978 m0 *1 0,71.76
X$978 61 62 63 221 64 222 257 258 cell_2rw
* cell instance $979 r0 *1 0,71.76
X$979 61 62 63 226 64 225 257 258 cell_2rw
* cell instance $980 m0 *1 0,74.75
X$980 61 62 63 231 64 232 257 258 cell_2rw
* cell instance $981 r0 *1 0,74.75
X$981 61 62 63 230 64 229 257 258 cell_2rw
* cell instance $982 m0 *1 0,77.74
X$982 61 62 63 227 64 228 257 258 cell_2rw
* cell instance $983 m0 *1 0,80.73
X$983 61 62 63 233 64 236 257 258 cell_2rw
* cell instance $984 r0 *1 0,77.74
X$984 61 62 63 237 64 238 257 258 cell_2rw
* cell instance $985 r0 *1 0,80.73
X$985 61 62 63 235 64 234 257 258 cell_2rw
* cell instance $986 m0 *1 0,83.72
X$986 61 62 63 240 64 242 257 258 cell_2rw
* cell instance $987 m0 *1 0,86.71
X$987 61 62 63 244 64 243 257 258 cell_2rw
* cell instance $988 r0 *1 0,83.72
X$988 61 62 63 239 64 241 257 258 cell_2rw
* cell instance $989 r0 *1 0,86.71
X$989 61 62 63 245 64 247 257 258 cell_2rw
* cell instance $990 m0 *1 0,89.7
X$990 61 62 63 250 64 249 257 258 cell_2rw
* cell instance $991 r0 *1 0,89.7
X$991 61 62 63 246 64 248 257 258 cell_2rw
* cell instance $992 m0 *1 0,92.69
X$992 61 62 63 253 64 256 257 258 cell_2rw
* cell instance $993 r0 *1 0,92.69
X$993 61 62 63 255 64 254 257 258 cell_2rw
* cell instance $994 m0 *1 0,95.68
X$994 61 62 63 251 64 252 257 258 cell_2rw
* cell instance $995 r0 *1 1.175,44.85
X$995 65 66 67 127 68 128 257 258 cell_2rw
* cell instance $996 m0 *1 1.175,47.84
X$996 65 66 67 126 68 125 257 258 cell_2rw
* cell instance $997 m0 *1 1.175,50.83
X$997 65 66 67 195 68 197 257 258 cell_2rw
* cell instance $998 r0 *1 1.175,47.84
X$998 65 66 67 199 68 201 257 258 cell_2rw
* cell instance $999 r0 *1 1.175,50.83
X$999 65 66 67 202 68 194 257 258 cell_2rw
* cell instance $1000 m0 *1 1.175,53.82
X$1000 65 66 67 198 68 193 257 258 cell_2rw
* cell instance $1001 r0 *1 1.175,53.82
X$1001 65 66 67 196 68 200 257 258 cell_2rw
* cell instance $1002 m0 *1 1.175,56.81
X$1002 65 66 67 203 68 207 257 258 cell_2rw
* cell instance $1003 r0 *1 1.175,56.81
X$1003 65 66 67 206 68 208 257 258 cell_2rw
* cell instance $1004 m0 *1 1.175,59.8
X$1004 65 66 67 205 68 204 257 258 cell_2rw
* cell instance $1005 r0 *1 1.175,59.8
X$1005 65 66 67 214 68 213 257 258 cell_2rw
* cell instance $1006 m0 *1 1.175,62.79
X$1006 65 66 67 212 68 211 257 258 cell_2rw
* cell instance $1007 r0 *1 1.175,62.79
X$1007 65 66 67 210 68 209 257 258 cell_2rw
* cell instance $1008 m0 *1 1.175,65.78
X$1008 65 66 67 219 68 217 257 258 cell_2rw
* cell instance $1009 r0 *1 1.175,65.78
X$1009 65 66 67 216 68 215 257 258 cell_2rw
* cell instance $1010 m0 *1 1.175,68.77
X$1010 65 66 67 218 68 220 257 258 cell_2rw
* cell instance $1011 r0 *1 1.175,68.77
X$1011 65 66 67 224 68 223 257 258 cell_2rw
* cell instance $1012 m0 *1 1.175,71.76
X$1012 65 66 67 221 68 222 257 258 cell_2rw
* cell instance $1013 r0 *1 1.175,71.76
X$1013 65 66 67 226 68 225 257 258 cell_2rw
* cell instance $1014 m0 *1 1.175,74.75
X$1014 65 66 67 231 68 232 257 258 cell_2rw
* cell instance $1015 r0 *1 1.175,74.75
X$1015 65 66 67 230 68 229 257 258 cell_2rw
* cell instance $1016 m0 *1 1.175,77.74
X$1016 65 66 67 227 68 228 257 258 cell_2rw
* cell instance $1017 r0 *1 1.175,77.74
X$1017 65 66 67 237 68 238 257 258 cell_2rw
* cell instance $1018 m0 *1 1.175,80.73
X$1018 65 66 67 233 68 236 257 258 cell_2rw
* cell instance $1019 m0 *1 1.175,83.72
X$1019 65 66 67 240 68 242 257 258 cell_2rw
* cell instance $1020 r0 *1 1.175,80.73
X$1020 65 66 67 235 68 234 257 258 cell_2rw
* cell instance $1021 r0 *1 1.175,83.72
X$1021 65 66 67 239 68 241 257 258 cell_2rw
* cell instance $1022 m0 *1 1.175,86.71
X$1022 65 66 67 244 68 243 257 258 cell_2rw
* cell instance $1023 r0 *1 1.175,86.71
X$1023 65 66 67 245 68 247 257 258 cell_2rw
* cell instance $1024 m0 *1 1.175,89.7
X$1024 65 66 67 250 68 249 257 258 cell_2rw
* cell instance $1025 r0 *1 1.175,89.7
X$1025 65 66 67 246 68 248 257 258 cell_2rw
* cell instance $1026 m0 *1 1.175,92.69
X$1026 65 66 67 253 68 256 257 258 cell_2rw
* cell instance $1027 r0 *1 1.175,92.69
X$1027 65 66 67 255 68 254 257 258 cell_2rw
* cell instance $1028 m0 *1 1.175,95.68
X$1028 65 66 67 251 68 252 257 258 cell_2rw
* cell instance $1029 m0 *1 2.35,47.84
X$1029 69 70 71 126 72 125 257 258 cell_2rw
* cell instance $1030 r0 *1 2.35,44.85
X$1030 69 70 71 127 72 128 257 258 cell_2rw
* cell instance $1031 r0 *1 2.35,47.84
X$1031 69 70 71 199 72 201 257 258 cell_2rw
* cell instance $1032 m0 *1 2.35,50.83
X$1032 69 70 71 195 72 197 257 258 cell_2rw
* cell instance $1033 r0 *1 2.35,50.83
X$1033 69 70 71 202 72 194 257 258 cell_2rw
* cell instance $1034 m0 *1 2.35,53.82
X$1034 69 70 71 198 72 193 257 258 cell_2rw
* cell instance $1035 m0 *1 2.35,56.81
X$1035 69 70 71 203 72 207 257 258 cell_2rw
* cell instance $1036 r0 *1 2.35,53.82
X$1036 69 70 71 196 72 200 257 258 cell_2rw
* cell instance $1037 r0 *1 2.35,56.81
X$1037 69 70 71 206 72 208 257 258 cell_2rw
* cell instance $1038 m0 *1 2.35,59.8
X$1038 69 70 71 205 72 204 257 258 cell_2rw
* cell instance $1039 m0 *1 2.35,62.79
X$1039 69 70 71 212 72 211 257 258 cell_2rw
* cell instance $1040 r0 *1 2.35,59.8
X$1040 69 70 71 214 72 213 257 258 cell_2rw
* cell instance $1041 r0 *1 2.35,62.79
X$1041 69 70 71 210 72 209 257 258 cell_2rw
* cell instance $1042 m0 *1 2.35,65.78
X$1042 69 70 71 219 72 217 257 258 cell_2rw
* cell instance $1043 r0 *1 2.35,65.78
X$1043 69 70 71 216 72 215 257 258 cell_2rw
* cell instance $1044 m0 *1 2.35,68.77
X$1044 69 70 71 218 72 220 257 258 cell_2rw
* cell instance $1045 m0 *1 2.35,71.76
X$1045 69 70 71 221 72 222 257 258 cell_2rw
* cell instance $1046 r0 *1 2.35,68.77
X$1046 69 70 71 224 72 223 257 258 cell_2rw
* cell instance $1047 m0 *1 2.35,74.75
X$1047 69 70 71 231 72 232 257 258 cell_2rw
* cell instance $1048 r0 *1 2.35,71.76
X$1048 69 70 71 226 72 225 257 258 cell_2rw
* cell instance $1049 r0 *1 2.35,74.75
X$1049 69 70 71 230 72 229 257 258 cell_2rw
* cell instance $1050 m0 *1 2.35,77.74
X$1050 69 70 71 227 72 228 257 258 cell_2rw
* cell instance $1051 r0 *1 2.35,77.74
X$1051 69 70 71 237 72 238 257 258 cell_2rw
* cell instance $1052 m0 *1 2.35,80.73
X$1052 69 70 71 233 72 236 257 258 cell_2rw
* cell instance $1053 r0 *1 2.35,80.73
X$1053 69 70 71 235 72 234 257 258 cell_2rw
* cell instance $1054 m0 *1 2.35,83.72
X$1054 69 70 71 240 72 242 257 258 cell_2rw
* cell instance $1055 m0 *1 2.35,86.71
X$1055 69 70 71 244 72 243 257 258 cell_2rw
* cell instance $1056 r0 *1 2.35,83.72
X$1056 69 70 71 239 72 241 257 258 cell_2rw
* cell instance $1057 r0 *1 2.35,86.71
X$1057 69 70 71 245 72 247 257 258 cell_2rw
* cell instance $1058 m0 *1 2.35,89.7
X$1058 69 70 71 250 72 249 257 258 cell_2rw
* cell instance $1059 r0 *1 2.35,89.7
X$1059 69 70 71 246 72 248 257 258 cell_2rw
* cell instance $1060 m0 *1 2.35,92.69
X$1060 69 70 71 253 72 256 257 258 cell_2rw
* cell instance $1061 r0 *1 2.35,92.69
X$1061 69 70 71 255 72 254 257 258 cell_2rw
* cell instance $1062 m0 *1 2.35,95.68
X$1062 69 70 71 251 72 252 257 258 cell_2rw
* cell instance $1063 r0 *1 3.525,44.85
X$1063 73 74 75 127 76 128 257 258 cell_2rw
* cell instance $1064 m0 *1 3.525,47.84
X$1064 73 74 75 126 76 125 257 258 cell_2rw
* cell instance $1065 m0 *1 3.525,50.83
X$1065 73 74 75 195 76 197 257 258 cell_2rw
* cell instance $1066 r0 *1 3.525,47.84
X$1066 73 74 75 199 76 201 257 258 cell_2rw
* cell instance $1067 r0 *1 3.525,50.83
X$1067 73 74 75 202 76 194 257 258 cell_2rw
* cell instance $1068 m0 *1 3.525,53.82
X$1068 73 74 75 198 76 193 257 258 cell_2rw
* cell instance $1069 r0 *1 3.525,53.82
X$1069 73 74 75 196 76 200 257 258 cell_2rw
* cell instance $1070 m0 *1 3.525,56.81
X$1070 73 74 75 203 76 207 257 258 cell_2rw
* cell instance $1071 m0 *1 3.525,59.8
X$1071 73 74 75 205 76 204 257 258 cell_2rw
* cell instance $1072 r0 *1 3.525,56.81
X$1072 73 74 75 206 76 208 257 258 cell_2rw
* cell instance $1073 r0 *1 3.525,59.8
X$1073 73 74 75 214 76 213 257 258 cell_2rw
* cell instance $1074 m0 *1 3.525,62.79
X$1074 73 74 75 212 76 211 257 258 cell_2rw
* cell instance $1075 r0 *1 3.525,62.79
X$1075 73 74 75 210 76 209 257 258 cell_2rw
* cell instance $1076 m0 *1 3.525,65.78
X$1076 73 74 75 219 76 217 257 258 cell_2rw
* cell instance $1077 r0 *1 3.525,65.78
X$1077 73 74 75 216 76 215 257 258 cell_2rw
* cell instance $1078 m0 *1 3.525,68.77
X$1078 73 74 75 218 76 220 257 258 cell_2rw
* cell instance $1079 r0 *1 3.525,68.77
X$1079 73 74 75 224 76 223 257 258 cell_2rw
* cell instance $1080 m0 *1 3.525,71.76
X$1080 73 74 75 221 76 222 257 258 cell_2rw
* cell instance $1081 r0 *1 3.525,71.76
X$1081 73 74 75 226 76 225 257 258 cell_2rw
* cell instance $1082 m0 *1 3.525,74.75
X$1082 73 74 75 231 76 232 257 258 cell_2rw
* cell instance $1083 m0 *1 3.525,77.74
X$1083 73 74 75 227 76 228 257 258 cell_2rw
* cell instance $1084 r0 *1 3.525,74.75
X$1084 73 74 75 230 76 229 257 258 cell_2rw
* cell instance $1085 r0 *1 3.525,77.74
X$1085 73 74 75 237 76 238 257 258 cell_2rw
* cell instance $1086 m0 *1 3.525,80.73
X$1086 73 74 75 233 76 236 257 258 cell_2rw
* cell instance $1087 r0 *1 3.525,80.73
X$1087 73 74 75 235 76 234 257 258 cell_2rw
* cell instance $1088 m0 *1 3.525,83.72
X$1088 73 74 75 240 76 242 257 258 cell_2rw
* cell instance $1089 r0 *1 3.525,83.72
X$1089 73 74 75 239 76 241 257 258 cell_2rw
* cell instance $1090 m0 *1 3.525,86.71
X$1090 73 74 75 244 76 243 257 258 cell_2rw
* cell instance $1091 r0 *1 3.525,86.71
X$1091 73 74 75 245 76 247 257 258 cell_2rw
* cell instance $1092 m0 *1 3.525,89.7
X$1092 73 74 75 250 76 249 257 258 cell_2rw
* cell instance $1093 r0 *1 3.525,89.7
X$1093 73 74 75 246 76 248 257 258 cell_2rw
* cell instance $1094 m0 *1 3.525,92.69
X$1094 73 74 75 253 76 256 257 258 cell_2rw
* cell instance $1095 r0 *1 3.525,92.69
X$1095 73 74 75 255 76 254 257 258 cell_2rw
* cell instance $1096 m0 *1 3.525,95.68
X$1096 73 74 75 251 76 252 257 258 cell_2rw
* cell instance $1097 r0 *1 4.7,44.85
X$1097 77 78 79 127 80 128 257 258 cell_2rw
* cell instance $1098 m0 *1 4.7,47.84
X$1098 77 78 79 126 80 125 257 258 cell_2rw
* cell instance $1099 r0 *1 4.7,47.84
X$1099 77 78 79 199 80 201 257 258 cell_2rw
* cell instance $1100 m0 *1 4.7,50.83
X$1100 77 78 79 195 80 197 257 258 cell_2rw
* cell instance $1101 r0 *1 4.7,50.83
X$1101 77 78 79 202 80 194 257 258 cell_2rw
* cell instance $1102 m0 *1 4.7,53.82
X$1102 77 78 79 198 80 193 257 258 cell_2rw
* cell instance $1103 r0 *1 4.7,53.82
X$1103 77 78 79 196 80 200 257 258 cell_2rw
* cell instance $1104 m0 *1 4.7,56.81
X$1104 77 78 79 203 80 207 257 258 cell_2rw
* cell instance $1105 r0 *1 4.7,56.81
X$1105 77 78 79 206 80 208 257 258 cell_2rw
* cell instance $1106 m0 *1 4.7,59.8
X$1106 77 78 79 205 80 204 257 258 cell_2rw
* cell instance $1107 r0 *1 4.7,59.8
X$1107 77 78 79 214 80 213 257 258 cell_2rw
* cell instance $1108 m0 *1 4.7,62.79
X$1108 77 78 79 212 80 211 257 258 cell_2rw
* cell instance $1109 r0 *1 4.7,62.79
X$1109 77 78 79 210 80 209 257 258 cell_2rw
* cell instance $1110 m0 *1 4.7,65.78
X$1110 77 78 79 219 80 217 257 258 cell_2rw
* cell instance $1111 m0 *1 4.7,68.77
X$1111 77 78 79 218 80 220 257 258 cell_2rw
* cell instance $1112 r0 *1 4.7,65.78
X$1112 77 78 79 216 80 215 257 258 cell_2rw
* cell instance $1113 r0 *1 4.7,68.77
X$1113 77 78 79 224 80 223 257 258 cell_2rw
* cell instance $1114 m0 *1 4.7,71.76
X$1114 77 78 79 221 80 222 257 258 cell_2rw
* cell instance $1115 m0 *1 4.7,74.75
X$1115 77 78 79 231 80 232 257 258 cell_2rw
* cell instance $1116 r0 *1 4.7,71.76
X$1116 77 78 79 226 80 225 257 258 cell_2rw
* cell instance $1117 r0 *1 4.7,74.75
X$1117 77 78 79 230 80 229 257 258 cell_2rw
* cell instance $1118 m0 *1 4.7,77.74
X$1118 77 78 79 227 80 228 257 258 cell_2rw
* cell instance $1119 r0 *1 4.7,77.74
X$1119 77 78 79 237 80 238 257 258 cell_2rw
* cell instance $1120 m0 *1 4.7,80.73
X$1120 77 78 79 233 80 236 257 258 cell_2rw
* cell instance $1121 r0 *1 4.7,80.73
X$1121 77 78 79 235 80 234 257 258 cell_2rw
* cell instance $1122 m0 *1 4.7,83.72
X$1122 77 78 79 240 80 242 257 258 cell_2rw
* cell instance $1123 m0 *1 4.7,86.71
X$1123 77 78 79 244 80 243 257 258 cell_2rw
* cell instance $1124 r0 *1 4.7,83.72
X$1124 77 78 79 239 80 241 257 258 cell_2rw
* cell instance $1125 m0 *1 4.7,89.7
X$1125 77 78 79 250 80 249 257 258 cell_2rw
* cell instance $1126 r0 *1 4.7,86.71
X$1126 77 78 79 245 80 247 257 258 cell_2rw
* cell instance $1127 r0 *1 4.7,89.7
X$1127 77 78 79 246 80 248 257 258 cell_2rw
* cell instance $1128 m0 *1 4.7,92.69
X$1128 77 78 79 253 80 256 257 258 cell_2rw
* cell instance $1129 r0 *1 4.7,92.69
X$1129 77 78 79 255 80 254 257 258 cell_2rw
* cell instance $1130 m0 *1 4.7,95.68
X$1130 77 78 79 251 80 252 257 258 cell_2rw
* cell instance $1131 m0 *1 5.875,47.84
X$1131 81 82 83 126 84 125 257 258 cell_2rw
* cell instance $1132 r0 *1 5.875,44.85
X$1132 81 82 83 127 84 128 257 258 cell_2rw
* cell instance $1133 r0 *1 5.875,47.84
X$1133 81 82 83 199 84 201 257 258 cell_2rw
* cell instance $1134 m0 *1 5.875,50.83
X$1134 81 82 83 195 84 197 257 258 cell_2rw
* cell instance $1135 r0 *1 5.875,50.83
X$1135 81 82 83 202 84 194 257 258 cell_2rw
* cell instance $1136 m0 *1 5.875,53.82
X$1136 81 82 83 198 84 193 257 258 cell_2rw
* cell instance $1137 r0 *1 5.875,53.82
X$1137 81 82 83 196 84 200 257 258 cell_2rw
* cell instance $1138 m0 *1 5.875,56.81
X$1138 81 82 83 203 84 207 257 258 cell_2rw
* cell instance $1139 r0 *1 5.875,56.81
X$1139 81 82 83 206 84 208 257 258 cell_2rw
* cell instance $1140 m0 *1 5.875,59.8
X$1140 81 82 83 205 84 204 257 258 cell_2rw
* cell instance $1141 r0 *1 5.875,59.8
X$1141 81 82 83 214 84 213 257 258 cell_2rw
* cell instance $1142 m0 *1 5.875,62.79
X$1142 81 82 83 212 84 211 257 258 cell_2rw
* cell instance $1143 r0 *1 5.875,62.79
X$1143 81 82 83 210 84 209 257 258 cell_2rw
* cell instance $1144 m0 *1 5.875,65.78
X$1144 81 82 83 219 84 217 257 258 cell_2rw
* cell instance $1145 r0 *1 5.875,65.78
X$1145 81 82 83 216 84 215 257 258 cell_2rw
* cell instance $1146 m0 *1 5.875,68.77
X$1146 81 82 83 218 84 220 257 258 cell_2rw
* cell instance $1147 r0 *1 5.875,68.77
X$1147 81 82 83 224 84 223 257 258 cell_2rw
* cell instance $1148 m0 *1 5.875,71.76
X$1148 81 82 83 221 84 222 257 258 cell_2rw
* cell instance $1149 r0 *1 5.875,71.76
X$1149 81 82 83 226 84 225 257 258 cell_2rw
* cell instance $1150 m0 *1 5.875,74.75
X$1150 81 82 83 231 84 232 257 258 cell_2rw
* cell instance $1151 m0 *1 5.875,77.74
X$1151 81 82 83 227 84 228 257 258 cell_2rw
* cell instance $1152 r0 *1 5.875,74.75
X$1152 81 82 83 230 84 229 257 258 cell_2rw
* cell instance $1153 r0 *1 5.875,77.74
X$1153 81 82 83 237 84 238 257 258 cell_2rw
* cell instance $1154 m0 *1 5.875,80.73
X$1154 81 82 83 233 84 236 257 258 cell_2rw
* cell instance $1155 r0 *1 5.875,80.73
X$1155 81 82 83 235 84 234 257 258 cell_2rw
* cell instance $1156 m0 *1 5.875,83.72
X$1156 81 82 83 240 84 242 257 258 cell_2rw
* cell instance $1157 r0 *1 5.875,83.72
X$1157 81 82 83 239 84 241 257 258 cell_2rw
* cell instance $1158 m0 *1 5.875,86.71
X$1158 81 82 83 244 84 243 257 258 cell_2rw
* cell instance $1159 r0 *1 5.875,86.71
X$1159 81 82 83 245 84 247 257 258 cell_2rw
* cell instance $1160 m0 *1 5.875,89.7
X$1160 81 82 83 250 84 249 257 258 cell_2rw
* cell instance $1161 r0 *1 5.875,89.7
X$1161 81 82 83 246 84 248 257 258 cell_2rw
* cell instance $1162 m0 *1 5.875,92.69
X$1162 81 82 83 253 84 256 257 258 cell_2rw
* cell instance $1163 r0 *1 5.875,92.69
X$1163 81 82 83 255 84 254 257 258 cell_2rw
* cell instance $1164 m0 *1 5.875,95.68
X$1164 81 82 83 251 84 252 257 258 cell_2rw
* cell instance $1165 r0 *1 7.05,44.85
X$1165 85 86 87 127 88 128 257 258 cell_2rw
* cell instance $1166 m0 *1 7.05,47.84
X$1166 85 86 87 126 88 125 257 258 cell_2rw
* cell instance $1167 r0 *1 7.05,47.84
X$1167 85 86 87 199 88 201 257 258 cell_2rw
* cell instance $1168 m0 *1 7.05,50.83
X$1168 85 86 87 195 88 197 257 258 cell_2rw
* cell instance $1169 r0 *1 7.05,50.83
X$1169 85 86 87 202 88 194 257 258 cell_2rw
* cell instance $1170 m0 *1 7.05,53.82
X$1170 85 86 87 198 88 193 257 258 cell_2rw
* cell instance $1171 r0 *1 7.05,53.82
X$1171 85 86 87 196 88 200 257 258 cell_2rw
* cell instance $1172 m0 *1 7.05,56.81
X$1172 85 86 87 203 88 207 257 258 cell_2rw
* cell instance $1173 r0 *1 7.05,56.81
X$1173 85 86 87 206 88 208 257 258 cell_2rw
* cell instance $1174 m0 *1 7.05,59.8
X$1174 85 86 87 205 88 204 257 258 cell_2rw
* cell instance $1175 r0 *1 7.05,59.8
X$1175 85 86 87 214 88 213 257 258 cell_2rw
* cell instance $1176 m0 *1 7.05,62.79
X$1176 85 86 87 212 88 211 257 258 cell_2rw
* cell instance $1177 r0 *1 7.05,62.79
X$1177 85 86 87 210 88 209 257 258 cell_2rw
* cell instance $1178 m0 *1 7.05,65.78
X$1178 85 86 87 219 88 217 257 258 cell_2rw
* cell instance $1179 r0 *1 7.05,65.78
X$1179 85 86 87 216 88 215 257 258 cell_2rw
* cell instance $1180 m0 *1 7.05,68.77
X$1180 85 86 87 218 88 220 257 258 cell_2rw
* cell instance $1181 r0 *1 7.05,68.77
X$1181 85 86 87 224 88 223 257 258 cell_2rw
* cell instance $1182 m0 *1 7.05,71.76
X$1182 85 86 87 221 88 222 257 258 cell_2rw
* cell instance $1183 r0 *1 7.05,71.76
X$1183 85 86 87 226 88 225 257 258 cell_2rw
* cell instance $1184 m0 *1 7.05,74.75
X$1184 85 86 87 231 88 232 257 258 cell_2rw
* cell instance $1185 r0 *1 7.05,74.75
X$1185 85 86 87 230 88 229 257 258 cell_2rw
* cell instance $1186 m0 *1 7.05,77.74
X$1186 85 86 87 227 88 228 257 258 cell_2rw
* cell instance $1187 r0 *1 7.05,77.74
X$1187 85 86 87 237 88 238 257 258 cell_2rw
* cell instance $1188 m0 *1 7.05,80.73
X$1188 85 86 87 233 88 236 257 258 cell_2rw
* cell instance $1189 m0 *1 7.05,83.72
X$1189 85 86 87 240 88 242 257 258 cell_2rw
* cell instance $1190 r0 *1 7.05,80.73
X$1190 85 86 87 235 88 234 257 258 cell_2rw
* cell instance $1191 r0 *1 7.05,83.72
X$1191 85 86 87 239 88 241 257 258 cell_2rw
* cell instance $1192 m0 *1 7.05,86.71
X$1192 85 86 87 244 88 243 257 258 cell_2rw
* cell instance $1193 r0 *1 7.05,86.71
X$1193 85 86 87 245 88 247 257 258 cell_2rw
* cell instance $1194 m0 *1 7.05,89.7
X$1194 85 86 87 250 88 249 257 258 cell_2rw
* cell instance $1195 m0 *1 7.05,92.69
X$1195 85 86 87 253 88 256 257 258 cell_2rw
* cell instance $1196 r0 *1 7.05,89.7
X$1196 85 86 87 246 88 248 257 258 cell_2rw
* cell instance $1197 m0 *1 7.05,95.68
X$1197 85 86 87 251 88 252 257 258 cell_2rw
* cell instance $1198 r0 *1 7.05,92.69
X$1198 85 86 87 255 88 254 257 258 cell_2rw
* cell instance $1199 m0 *1 8.225,47.84
X$1199 89 90 91 126 92 125 257 258 cell_2rw
* cell instance $1200 r0 *1 8.225,44.85
X$1200 89 90 91 127 92 128 257 258 cell_2rw
* cell instance $1201 m0 *1 8.225,50.83
X$1201 89 90 91 195 92 197 257 258 cell_2rw
* cell instance $1202 r0 *1 8.225,47.84
X$1202 89 90 91 199 92 201 257 258 cell_2rw
* cell instance $1203 r0 *1 8.225,50.83
X$1203 89 90 91 202 92 194 257 258 cell_2rw
* cell instance $1204 m0 *1 8.225,53.82
X$1204 89 90 91 198 92 193 257 258 cell_2rw
* cell instance $1205 r0 *1 8.225,53.82
X$1205 89 90 91 196 92 200 257 258 cell_2rw
* cell instance $1206 m0 *1 8.225,56.81
X$1206 89 90 91 203 92 207 257 258 cell_2rw
* cell instance $1207 r0 *1 8.225,56.81
X$1207 89 90 91 206 92 208 257 258 cell_2rw
* cell instance $1208 m0 *1 8.225,59.8
X$1208 89 90 91 205 92 204 257 258 cell_2rw
* cell instance $1209 r0 *1 8.225,59.8
X$1209 89 90 91 214 92 213 257 258 cell_2rw
* cell instance $1210 m0 *1 8.225,62.79
X$1210 89 90 91 212 92 211 257 258 cell_2rw
* cell instance $1211 r0 *1 8.225,62.79
X$1211 89 90 91 210 92 209 257 258 cell_2rw
* cell instance $1212 m0 *1 8.225,65.78
X$1212 89 90 91 219 92 217 257 258 cell_2rw
* cell instance $1213 r0 *1 8.225,65.78
X$1213 89 90 91 216 92 215 257 258 cell_2rw
* cell instance $1214 m0 *1 8.225,68.77
X$1214 89 90 91 218 92 220 257 258 cell_2rw
* cell instance $1215 m0 *1 8.225,71.76
X$1215 89 90 91 221 92 222 257 258 cell_2rw
* cell instance $1216 r0 *1 8.225,68.77
X$1216 89 90 91 224 92 223 257 258 cell_2rw
* cell instance $1217 m0 *1 8.225,74.75
X$1217 89 90 91 231 92 232 257 258 cell_2rw
* cell instance $1218 r0 *1 8.225,71.76
X$1218 89 90 91 226 92 225 257 258 cell_2rw
* cell instance $1219 r0 *1 8.225,74.75
X$1219 89 90 91 230 92 229 257 258 cell_2rw
* cell instance $1220 m0 *1 8.225,77.74
X$1220 89 90 91 227 92 228 257 258 cell_2rw
* cell instance $1221 r0 *1 8.225,77.74
X$1221 89 90 91 237 92 238 257 258 cell_2rw
* cell instance $1222 m0 *1 8.225,80.73
X$1222 89 90 91 233 92 236 257 258 cell_2rw
* cell instance $1223 r0 *1 8.225,80.73
X$1223 89 90 91 235 92 234 257 258 cell_2rw
* cell instance $1224 m0 *1 8.225,83.72
X$1224 89 90 91 240 92 242 257 258 cell_2rw
* cell instance $1225 r0 *1 8.225,83.72
X$1225 89 90 91 239 92 241 257 258 cell_2rw
* cell instance $1226 m0 *1 8.225,86.71
X$1226 89 90 91 244 92 243 257 258 cell_2rw
* cell instance $1227 r0 *1 8.225,86.71
X$1227 89 90 91 245 92 247 257 258 cell_2rw
* cell instance $1228 m0 *1 8.225,89.7
X$1228 89 90 91 250 92 249 257 258 cell_2rw
* cell instance $1229 r0 *1 8.225,89.7
X$1229 89 90 91 246 92 248 257 258 cell_2rw
* cell instance $1230 m0 *1 8.225,92.69
X$1230 89 90 91 253 92 256 257 258 cell_2rw
* cell instance $1231 m0 *1 8.225,95.68
X$1231 89 90 91 251 92 252 257 258 cell_2rw
* cell instance $1232 r0 *1 8.225,92.69
X$1232 89 90 91 255 92 254 257 258 cell_2rw
* cell instance $1233 r0 *1 9.4,44.85
X$1233 93 94 95 127 96 128 257 258 cell_2rw
* cell instance $1234 m0 *1 9.4,47.84
X$1234 93 94 95 126 96 125 257 258 cell_2rw
* cell instance $1235 r0 *1 9.4,47.84
X$1235 93 94 95 199 96 201 257 258 cell_2rw
* cell instance $1236 m0 *1 9.4,50.83
X$1236 93 94 95 195 96 197 257 258 cell_2rw
* cell instance $1237 r0 *1 9.4,50.83
X$1237 93 94 95 202 96 194 257 258 cell_2rw
* cell instance $1238 m0 *1 9.4,53.82
X$1238 93 94 95 198 96 193 257 258 cell_2rw
* cell instance $1239 r0 *1 9.4,53.82
X$1239 93 94 95 196 96 200 257 258 cell_2rw
* cell instance $1240 m0 *1 9.4,56.81
X$1240 93 94 95 203 96 207 257 258 cell_2rw
* cell instance $1241 r0 *1 9.4,56.81
X$1241 93 94 95 206 96 208 257 258 cell_2rw
* cell instance $1242 m0 *1 9.4,59.8
X$1242 93 94 95 205 96 204 257 258 cell_2rw
* cell instance $1243 m0 *1 9.4,62.79
X$1243 93 94 95 212 96 211 257 258 cell_2rw
* cell instance $1244 r0 *1 9.4,59.8
X$1244 93 94 95 214 96 213 257 258 cell_2rw
* cell instance $1245 r0 *1 9.4,62.79
X$1245 93 94 95 210 96 209 257 258 cell_2rw
* cell instance $1246 m0 *1 9.4,65.78
X$1246 93 94 95 219 96 217 257 258 cell_2rw
* cell instance $1247 r0 *1 9.4,65.78
X$1247 93 94 95 216 96 215 257 258 cell_2rw
* cell instance $1248 m0 *1 9.4,68.77
X$1248 93 94 95 218 96 220 257 258 cell_2rw
* cell instance $1249 r0 *1 9.4,68.77
X$1249 93 94 95 224 96 223 257 258 cell_2rw
* cell instance $1250 m0 *1 9.4,71.76
X$1250 93 94 95 221 96 222 257 258 cell_2rw
* cell instance $1251 r0 *1 9.4,71.76
X$1251 93 94 95 226 96 225 257 258 cell_2rw
* cell instance $1252 m0 *1 9.4,74.75
X$1252 93 94 95 231 96 232 257 258 cell_2rw
* cell instance $1253 r0 *1 9.4,74.75
X$1253 93 94 95 230 96 229 257 258 cell_2rw
* cell instance $1254 m0 *1 9.4,77.74
X$1254 93 94 95 227 96 228 257 258 cell_2rw
* cell instance $1255 r0 *1 9.4,77.74
X$1255 93 94 95 237 96 238 257 258 cell_2rw
* cell instance $1256 m0 *1 9.4,80.73
X$1256 93 94 95 233 96 236 257 258 cell_2rw
* cell instance $1257 r0 *1 9.4,80.73
X$1257 93 94 95 235 96 234 257 258 cell_2rw
* cell instance $1258 m0 *1 9.4,83.72
X$1258 93 94 95 240 96 242 257 258 cell_2rw
* cell instance $1259 r0 *1 9.4,83.72
X$1259 93 94 95 239 96 241 257 258 cell_2rw
* cell instance $1260 m0 *1 9.4,86.71
X$1260 93 94 95 244 96 243 257 258 cell_2rw
* cell instance $1261 m0 *1 9.4,89.7
X$1261 93 94 95 250 96 249 257 258 cell_2rw
* cell instance $1262 r0 *1 9.4,86.71
X$1262 93 94 95 245 96 247 257 258 cell_2rw
* cell instance $1263 r0 *1 9.4,89.7
X$1263 93 94 95 246 96 248 257 258 cell_2rw
* cell instance $1264 m0 *1 9.4,92.69
X$1264 93 94 95 253 96 256 257 258 cell_2rw
* cell instance $1265 m0 *1 9.4,95.68
X$1265 93 94 95 251 96 252 257 258 cell_2rw
* cell instance $1266 r0 *1 9.4,92.69
X$1266 93 94 95 255 96 254 257 258 cell_2rw
* cell instance $1267 r0 *1 10.575,44.85
X$1267 97 98 99 127 100 128 257 258 cell_2rw
* cell instance $1268 m0 *1 10.575,47.84
X$1268 97 98 99 126 100 125 257 258 cell_2rw
* cell instance $1269 r0 *1 10.575,47.84
X$1269 97 98 99 199 100 201 257 258 cell_2rw
* cell instance $1270 m0 *1 10.575,50.83
X$1270 97 98 99 195 100 197 257 258 cell_2rw
* cell instance $1271 r0 *1 10.575,50.83
X$1271 97 98 99 202 100 194 257 258 cell_2rw
* cell instance $1272 m0 *1 10.575,53.82
X$1272 97 98 99 198 100 193 257 258 cell_2rw
* cell instance $1273 r0 *1 10.575,53.82
X$1273 97 98 99 196 100 200 257 258 cell_2rw
* cell instance $1274 m0 *1 10.575,56.81
X$1274 97 98 99 203 100 207 257 258 cell_2rw
* cell instance $1275 r0 *1 10.575,56.81
X$1275 97 98 99 206 100 208 257 258 cell_2rw
* cell instance $1276 m0 *1 10.575,59.8
X$1276 97 98 99 205 100 204 257 258 cell_2rw
* cell instance $1277 r0 *1 10.575,59.8
X$1277 97 98 99 214 100 213 257 258 cell_2rw
* cell instance $1278 m0 *1 10.575,62.79
X$1278 97 98 99 212 100 211 257 258 cell_2rw
* cell instance $1279 r0 *1 10.575,62.79
X$1279 97 98 99 210 100 209 257 258 cell_2rw
* cell instance $1280 m0 *1 10.575,65.78
X$1280 97 98 99 219 100 217 257 258 cell_2rw
* cell instance $1281 r0 *1 10.575,65.78
X$1281 97 98 99 216 100 215 257 258 cell_2rw
* cell instance $1282 m0 *1 10.575,68.77
X$1282 97 98 99 218 100 220 257 258 cell_2rw
* cell instance $1283 r0 *1 10.575,68.77
X$1283 97 98 99 224 100 223 257 258 cell_2rw
* cell instance $1284 m0 *1 10.575,71.76
X$1284 97 98 99 221 100 222 257 258 cell_2rw
* cell instance $1285 r0 *1 10.575,71.76
X$1285 97 98 99 226 100 225 257 258 cell_2rw
* cell instance $1286 m0 *1 10.575,74.75
X$1286 97 98 99 231 100 232 257 258 cell_2rw
* cell instance $1287 r0 *1 10.575,74.75
X$1287 97 98 99 230 100 229 257 258 cell_2rw
* cell instance $1288 m0 *1 10.575,77.74
X$1288 97 98 99 227 100 228 257 258 cell_2rw
* cell instance $1289 r0 *1 10.575,77.74
X$1289 97 98 99 237 100 238 257 258 cell_2rw
* cell instance $1290 m0 *1 10.575,80.73
X$1290 97 98 99 233 100 236 257 258 cell_2rw
* cell instance $1291 r0 *1 10.575,80.73
X$1291 97 98 99 235 100 234 257 258 cell_2rw
* cell instance $1292 m0 *1 10.575,83.72
X$1292 97 98 99 240 100 242 257 258 cell_2rw
* cell instance $1293 m0 *1 10.575,86.71
X$1293 97 98 99 244 100 243 257 258 cell_2rw
* cell instance $1294 r0 *1 10.575,83.72
X$1294 97 98 99 239 100 241 257 258 cell_2rw
* cell instance $1295 r0 *1 10.575,86.71
X$1295 97 98 99 245 100 247 257 258 cell_2rw
* cell instance $1296 m0 *1 10.575,89.7
X$1296 97 98 99 250 100 249 257 258 cell_2rw
* cell instance $1297 r0 *1 10.575,89.7
X$1297 97 98 99 246 100 248 257 258 cell_2rw
* cell instance $1298 m0 *1 10.575,92.69
X$1298 97 98 99 253 100 256 257 258 cell_2rw
* cell instance $1299 m0 *1 10.575,95.68
X$1299 97 98 99 251 100 252 257 258 cell_2rw
* cell instance $1300 r0 *1 10.575,92.69
X$1300 97 98 99 255 100 254 257 258 cell_2rw
* cell instance $1301 m0 *1 11.75,47.84
X$1301 101 102 103 126 104 125 257 258 cell_2rw
* cell instance $1302 r0 *1 11.75,44.85
X$1302 101 102 103 127 104 128 257 258 cell_2rw
* cell instance $1303 r0 *1 11.75,47.84
X$1303 101 102 103 199 104 201 257 258 cell_2rw
* cell instance $1304 m0 *1 11.75,50.83
X$1304 101 102 103 195 104 197 257 258 cell_2rw
* cell instance $1305 m0 *1 11.75,53.82
X$1305 101 102 103 198 104 193 257 258 cell_2rw
* cell instance $1306 r0 *1 11.75,50.83
X$1306 101 102 103 202 104 194 257 258 cell_2rw
* cell instance $1307 r0 *1 11.75,53.82
X$1307 101 102 103 196 104 200 257 258 cell_2rw
* cell instance $1308 m0 *1 11.75,56.81
X$1308 101 102 103 203 104 207 257 258 cell_2rw
* cell instance $1309 r0 *1 11.75,56.81
X$1309 101 102 103 206 104 208 257 258 cell_2rw
* cell instance $1310 m0 *1 11.75,59.8
X$1310 101 102 103 205 104 204 257 258 cell_2rw
* cell instance $1311 r0 *1 11.75,59.8
X$1311 101 102 103 214 104 213 257 258 cell_2rw
* cell instance $1312 m0 *1 11.75,62.79
X$1312 101 102 103 212 104 211 257 258 cell_2rw
* cell instance $1313 m0 *1 11.75,65.78
X$1313 101 102 103 219 104 217 257 258 cell_2rw
* cell instance $1314 r0 *1 11.75,62.79
X$1314 101 102 103 210 104 209 257 258 cell_2rw
* cell instance $1315 m0 *1 11.75,68.77
X$1315 101 102 103 218 104 220 257 258 cell_2rw
* cell instance $1316 r0 *1 11.75,65.78
X$1316 101 102 103 216 104 215 257 258 cell_2rw
* cell instance $1317 r0 *1 11.75,68.77
X$1317 101 102 103 224 104 223 257 258 cell_2rw
* cell instance $1318 m0 *1 11.75,71.76
X$1318 101 102 103 221 104 222 257 258 cell_2rw
* cell instance $1319 r0 *1 11.75,71.76
X$1319 101 102 103 226 104 225 257 258 cell_2rw
* cell instance $1320 m0 *1 11.75,74.75
X$1320 101 102 103 231 104 232 257 258 cell_2rw
* cell instance $1321 r0 *1 11.75,74.75
X$1321 101 102 103 230 104 229 257 258 cell_2rw
* cell instance $1322 m0 *1 11.75,77.74
X$1322 101 102 103 227 104 228 257 258 cell_2rw
* cell instance $1323 r0 *1 11.75,77.74
X$1323 101 102 103 237 104 238 257 258 cell_2rw
* cell instance $1324 m0 *1 11.75,80.73
X$1324 101 102 103 233 104 236 257 258 cell_2rw
* cell instance $1325 r0 *1 11.75,80.73
X$1325 101 102 103 235 104 234 257 258 cell_2rw
* cell instance $1326 m0 *1 11.75,83.72
X$1326 101 102 103 240 104 242 257 258 cell_2rw
* cell instance $1327 m0 *1 11.75,86.71
X$1327 101 102 103 244 104 243 257 258 cell_2rw
* cell instance $1328 r0 *1 11.75,83.72
X$1328 101 102 103 239 104 241 257 258 cell_2rw
* cell instance $1329 r0 *1 11.75,86.71
X$1329 101 102 103 245 104 247 257 258 cell_2rw
* cell instance $1330 m0 *1 11.75,89.7
X$1330 101 102 103 250 104 249 257 258 cell_2rw
* cell instance $1331 r0 *1 11.75,89.7
X$1331 101 102 103 246 104 248 257 258 cell_2rw
* cell instance $1332 m0 *1 11.75,92.69
X$1332 101 102 103 253 104 256 257 258 cell_2rw
* cell instance $1333 r0 *1 11.75,92.69
X$1333 101 102 103 255 104 254 257 258 cell_2rw
* cell instance $1334 m0 *1 11.75,95.68
X$1334 101 102 103 251 104 252 257 258 cell_2rw
* cell instance $1335 r0 *1 12.925,44.85
X$1335 105 106 107 127 108 128 257 258 cell_2rw
* cell instance $1336 m0 *1 12.925,47.84
X$1336 105 106 107 126 108 125 257 258 cell_2rw
* cell instance $1337 m0 *1 12.925,50.83
X$1337 105 106 107 195 108 197 257 258 cell_2rw
* cell instance $1338 r0 *1 12.925,47.84
X$1338 105 106 107 199 108 201 257 258 cell_2rw
* cell instance $1339 m0 *1 12.925,53.82
X$1339 105 106 107 198 108 193 257 258 cell_2rw
* cell instance $1340 r0 *1 12.925,50.83
X$1340 105 106 107 202 108 194 257 258 cell_2rw
* cell instance $1341 r0 *1 12.925,53.82
X$1341 105 106 107 196 108 200 257 258 cell_2rw
* cell instance $1342 m0 *1 12.925,56.81
X$1342 105 106 107 203 108 207 257 258 cell_2rw
* cell instance $1343 r0 *1 12.925,56.81
X$1343 105 106 107 206 108 208 257 258 cell_2rw
* cell instance $1344 m0 *1 12.925,59.8
X$1344 105 106 107 205 108 204 257 258 cell_2rw
* cell instance $1345 r0 *1 12.925,59.8
X$1345 105 106 107 214 108 213 257 258 cell_2rw
* cell instance $1346 m0 *1 12.925,62.79
X$1346 105 106 107 212 108 211 257 258 cell_2rw
* cell instance $1347 r0 *1 12.925,62.79
X$1347 105 106 107 210 108 209 257 258 cell_2rw
* cell instance $1348 m0 *1 12.925,65.78
X$1348 105 106 107 219 108 217 257 258 cell_2rw
* cell instance $1349 r0 *1 12.925,65.78
X$1349 105 106 107 216 108 215 257 258 cell_2rw
* cell instance $1350 m0 *1 12.925,68.77
X$1350 105 106 107 218 108 220 257 258 cell_2rw
* cell instance $1351 r0 *1 12.925,68.77
X$1351 105 106 107 224 108 223 257 258 cell_2rw
* cell instance $1352 m0 *1 12.925,71.76
X$1352 105 106 107 221 108 222 257 258 cell_2rw
* cell instance $1353 r0 *1 12.925,71.76
X$1353 105 106 107 226 108 225 257 258 cell_2rw
* cell instance $1354 m0 *1 12.925,74.75
X$1354 105 106 107 231 108 232 257 258 cell_2rw
* cell instance $1355 r0 *1 12.925,74.75
X$1355 105 106 107 230 108 229 257 258 cell_2rw
* cell instance $1356 m0 *1 12.925,77.74
X$1356 105 106 107 227 108 228 257 258 cell_2rw
* cell instance $1357 r0 *1 12.925,77.74
X$1357 105 106 107 237 108 238 257 258 cell_2rw
* cell instance $1358 m0 *1 12.925,80.73
X$1358 105 106 107 233 108 236 257 258 cell_2rw
* cell instance $1359 r0 *1 12.925,80.73
X$1359 105 106 107 235 108 234 257 258 cell_2rw
* cell instance $1360 m0 *1 12.925,83.72
X$1360 105 106 107 240 108 242 257 258 cell_2rw
* cell instance $1361 r0 *1 12.925,83.72
X$1361 105 106 107 239 108 241 257 258 cell_2rw
* cell instance $1362 m0 *1 12.925,86.71
X$1362 105 106 107 244 108 243 257 258 cell_2rw
* cell instance $1363 r0 *1 12.925,86.71
X$1363 105 106 107 245 108 247 257 258 cell_2rw
* cell instance $1364 m0 *1 12.925,89.7
X$1364 105 106 107 250 108 249 257 258 cell_2rw
* cell instance $1365 r0 *1 12.925,89.7
X$1365 105 106 107 246 108 248 257 258 cell_2rw
* cell instance $1366 m0 *1 12.925,92.69
X$1366 105 106 107 253 108 256 257 258 cell_2rw
* cell instance $1367 r0 *1 12.925,92.69
X$1367 105 106 107 255 108 254 257 258 cell_2rw
* cell instance $1368 m0 *1 12.925,95.68
X$1368 105 106 107 251 108 252 257 258 cell_2rw
* cell instance $1369 r0 *1 14.1,44.85
X$1369 109 110 111 127 112 128 257 258 cell_2rw
* cell instance $1370 m0 *1 14.1,47.84
X$1370 109 110 111 126 112 125 257 258 cell_2rw
* cell instance $1371 r0 *1 14.1,47.84
X$1371 109 110 111 199 112 201 257 258 cell_2rw
* cell instance $1372 m0 *1 14.1,50.83
X$1372 109 110 111 195 112 197 257 258 cell_2rw
* cell instance $1373 r0 *1 14.1,50.83
X$1373 109 110 111 202 112 194 257 258 cell_2rw
* cell instance $1374 m0 *1 14.1,53.82
X$1374 109 110 111 198 112 193 257 258 cell_2rw
* cell instance $1375 r0 *1 14.1,53.82
X$1375 109 110 111 196 112 200 257 258 cell_2rw
* cell instance $1376 m0 *1 14.1,56.81
X$1376 109 110 111 203 112 207 257 258 cell_2rw
* cell instance $1377 r0 *1 14.1,56.81
X$1377 109 110 111 206 112 208 257 258 cell_2rw
* cell instance $1378 m0 *1 14.1,59.8
X$1378 109 110 111 205 112 204 257 258 cell_2rw
* cell instance $1379 m0 *1 14.1,62.79
X$1379 109 110 111 212 112 211 257 258 cell_2rw
* cell instance $1380 r0 *1 14.1,59.8
X$1380 109 110 111 214 112 213 257 258 cell_2rw
* cell instance $1381 r0 *1 14.1,62.79
X$1381 109 110 111 210 112 209 257 258 cell_2rw
* cell instance $1382 m0 *1 14.1,65.78
X$1382 109 110 111 219 112 217 257 258 cell_2rw
* cell instance $1383 r0 *1 14.1,65.78
X$1383 109 110 111 216 112 215 257 258 cell_2rw
* cell instance $1384 m0 *1 14.1,68.77
X$1384 109 110 111 218 112 220 257 258 cell_2rw
* cell instance $1385 r0 *1 14.1,68.77
X$1385 109 110 111 224 112 223 257 258 cell_2rw
* cell instance $1386 m0 *1 14.1,71.76
X$1386 109 110 111 221 112 222 257 258 cell_2rw
* cell instance $1387 r0 *1 14.1,71.76
X$1387 109 110 111 226 112 225 257 258 cell_2rw
* cell instance $1388 m0 *1 14.1,74.75
X$1388 109 110 111 231 112 232 257 258 cell_2rw
* cell instance $1389 r0 *1 14.1,74.75
X$1389 109 110 111 230 112 229 257 258 cell_2rw
* cell instance $1390 m0 *1 14.1,77.74
X$1390 109 110 111 227 112 228 257 258 cell_2rw
* cell instance $1391 r0 *1 14.1,77.74
X$1391 109 110 111 237 112 238 257 258 cell_2rw
* cell instance $1392 m0 *1 14.1,80.73
X$1392 109 110 111 233 112 236 257 258 cell_2rw
* cell instance $1393 r0 *1 14.1,80.73
X$1393 109 110 111 235 112 234 257 258 cell_2rw
* cell instance $1394 m0 *1 14.1,83.72
X$1394 109 110 111 240 112 242 257 258 cell_2rw
* cell instance $1395 m0 *1 14.1,86.71
X$1395 109 110 111 244 112 243 257 258 cell_2rw
* cell instance $1396 r0 *1 14.1,83.72
X$1396 109 110 111 239 112 241 257 258 cell_2rw
* cell instance $1397 r0 *1 14.1,86.71
X$1397 109 110 111 245 112 247 257 258 cell_2rw
* cell instance $1398 m0 *1 14.1,89.7
X$1398 109 110 111 250 112 249 257 258 cell_2rw
* cell instance $1399 r0 *1 14.1,89.7
X$1399 109 110 111 246 112 248 257 258 cell_2rw
* cell instance $1400 m0 *1 14.1,92.69
X$1400 109 110 111 253 112 256 257 258 cell_2rw
* cell instance $1401 r0 *1 14.1,92.69
X$1401 109 110 111 255 112 254 257 258 cell_2rw
* cell instance $1402 m0 *1 14.1,95.68
X$1402 109 110 111 251 112 252 257 258 cell_2rw
* cell instance $1403 r0 *1 15.275,44.85
X$1403 113 114 115 127 116 128 257 258 cell_2rw
* cell instance $1404 m0 *1 15.275,47.84
X$1404 113 114 115 126 116 125 257 258 cell_2rw
* cell instance $1405 m0 *1 15.275,50.83
X$1405 113 114 115 195 116 197 257 258 cell_2rw
* cell instance $1406 r0 *1 15.275,47.84
X$1406 113 114 115 199 116 201 257 258 cell_2rw
* cell instance $1407 m0 *1 15.275,53.82
X$1407 113 114 115 198 116 193 257 258 cell_2rw
* cell instance $1408 r0 *1 15.275,50.83
X$1408 113 114 115 202 116 194 257 258 cell_2rw
* cell instance $1409 r0 *1 15.275,53.82
X$1409 113 114 115 196 116 200 257 258 cell_2rw
* cell instance $1410 m0 *1 15.275,56.81
X$1410 113 114 115 203 116 207 257 258 cell_2rw
* cell instance $1411 r0 *1 15.275,56.81
X$1411 113 114 115 206 116 208 257 258 cell_2rw
* cell instance $1412 m0 *1 15.275,59.8
X$1412 113 114 115 205 116 204 257 258 cell_2rw
* cell instance $1413 r0 *1 15.275,59.8
X$1413 113 114 115 214 116 213 257 258 cell_2rw
* cell instance $1414 m0 *1 15.275,62.79
X$1414 113 114 115 212 116 211 257 258 cell_2rw
* cell instance $1415 r0 *1 15.275,62.79
X$1415 113 114 115 210 116 209 257 258 cell_2rw
* cell instance $1416 m0 *1 15.275,65.78
X$1416 113 114 115 219 116 217 257 258 cell_2rw
* cell instance $1417 r0 *1 15.275,65.78
X$1417 113 114 115 216 116 215 257 258 cell_2rw
* cell instance $1418 m0 *1 15.275,68.77
X$1418 113 114 115 218 116 220 257 258 cell_2rw
* cell instance $1419 r0 *1 15.275,68.77
X$1419 113 114 115 224 116 223 257 258 cell_2rw
* cell instance $1420 m0 *1 15.275,71.76
X$1420 113 114 115 221 116 222 257 258 cell_2rw
* cell instance $1421 r0 *1 15.275,71.76
X$1421 113 114 115 226 116 225 257 258 cell_2rw
* cell instance $1422 m0 *1 15.275,74.75
X$1422 113 114 115 231 116 232 257 258 cell_2rw
* cell instance $1423 r0 *1 15.275,74.75
X$1423 113 114 115 230 116 229 257 258 cell_2rw
* cell instance $1424 m0 *1 15.275,77.74
X$1424 113 114 115 227 116 228 257 258 cell_2rw
* cell instance $1425 m0 *1 15.275,80.73
X$1425 113 114 115 233 116 236 257 258 cell_2rw
* cell instance $1426 r0 *1 15.275,77.74
X$1426 113 114 115 237 116 238 257 258 cell_2rw
* cell instance $1427 m0 *1 15.275,83.72
X$1427 113 114 115 240 116 242 257 258 cell_2rw
* cell instance $1428 r0 *1 15.275,80.73
X$1428 113 114 115 235 116 234 257 258 cell_2rw
* cell instance $1429 r0 *1 15.275,83.72
X$1429 113 114 115 239 116 241 257 258 cell_2rw
* cell instance $1430 m0 *1 15.275,86.71
X$1430 113 114 115 244 116 243 257 258 cell_2rw
* cell instance $1431 m0 *1 15.275,89.7
X$1431 113 114 115 250 116 249 257 258 cell_2rw
* cell instance $1432 r0 *1 15.275,86.71
X$1432 113 114 115 245 116 247 257 258 cell_2rw
* cell instance $1433 r0 *1 15.275,89.7
X$1433 113 114 115 246 116 248 257 258 cell_2rw
* cell instance $1434 m0 *1 15.275,92.69
X$1434 113 114 115 253 116 256 257 258 cell_2rw
* cell instance $1435 r0 *1 15.275,92.69
X$1435 113 114 115 255 116 254 257 258 cell_2rw
* cell instance $1436 m0 *1 15.275,95.68
X$1436 113 114 115 251 116 252 257 258 cell_2rw
* cell instance $1437 r0 *1 16.45,44.85
X$1437 117 118 119 127 120 128 257 258 cell_2rw
* cell instance $1438 m0 *1 16.45,47.84
X$1438 117 118 119 126 120 125 257 258 cell_2rw
* cell instance $1439 r0 *1 16.45,47.84
X$1439 117 118 119 199 120 201 257 258 cell_2rw
* cell instance $1440 m0 *1 16.45,50.83
X$1440 117 118 119 195 120 197 257 258 cell_2rw
* cell instance $1441 m0 *1 16.45,53.82
X$1441 117 118 119 198 120 193 257 258 cell_2rw
* cell instance $1442 r0 *1 16.45,50.83
X$1442 117 118 119 202 120 194 257 258 cell_2rw
* cell instance $1443 r0 *1 16.45,53.82
X$1443 117 118 119 196 120 200 257 258 cell_2rw
* cell instance $1444 m0 *1 16.45,56.81
X$1444 117 118 119 203 120 207 257 258 cell_2rw
* cell instance $1445 m0 *1 16.45,59.8
X$1445 117 118 119 205 120 204 257 258 cell_2rw
* cell instance $1446 r0 *1 16.45,56.81
X$1446 117 118 119 206 120 208 257 258 cell_2rw
* cell instance $1447 m0 *1 16.45,62.79
X$1447 117 118 119 212 120 211 257 258 cell_2rw
* cell instance $1448 r0 *1 16.45,59.8
X$1448 117 118 119 214 120 213 257 258 cell_2rw
* cell instance $1449 r0 *1 16.45,62.79
X$1449 117 118 119 210 120 209 257 258 cell_2rw
* cell instance $1450 m0 *1 16.45,65.78
X$1450 117 118 119 219 120 217 257 258 cell_2rw
* cell instance $1451 r0 *1 16.45,65.78
X$1451 117 118 119 216 120 215 257 258 cell_2rw
* cell instance $1452 m0 *1 16.45,68.77
X$1452 117 118 119 218 120 220 257 258 cell_2rw
* cell instance $1453 r0 *1 16.45,68.77
X$1453 117 118 119 224 120 223 257 258 cell_2rw
* cell instance $1454 m0 *1 16.45,71.76
X$1454 117 118 119 221 120 222 257 258 cell_2rw
* cell instance $1455 r0 *1 16.45,71.76
X$1455 117 118 119 226 120 225 257 258 cell_2rw
* cell instance $1456 m0 *1 16.45,74.75
X$1456 117 118 119 231 120 232 257 258 cell_2rw
* cell instance $1457 r0 *1 16.45,74.75
X$1457 117 118 119 230 120 229 257 258 cell_2rw
* cell instance $1458 m0 *1 16.45,77.74
X$1458 117 118 119 227 120 228 257 258 cell_2rw
* cell instance $1459 m0 *1 16.45,80.73
X$1459 117 118 119 233 120 236 257 258 cell_2rw
* cell instance $1460 r0 *1 16.45,77.74
X$1460 117 118 119 237 120 238 257 258 cell_2rw
* cell instance $1461 r0 *1 16.45,80.73
X$1461 117 118 119 235 120 234 257 258 cell_2rw
* cell instance $1462 m0 *1 16.45,83.72
X$1462 117 118 119 240 120 242 257 258 cell_2rw
* cell instance $1463 r0 *1 16.45,83.72
X$1463 117 118 119 239 120 241 257 258 cell_2rw
* cell instance $1464 m0 *1 16.45,86.71
X$1464 117 118 119 244 120 243 257 258 cell_2rw
* cell instance $1465 r0 *1 16.45,86.71
X$1465 117 118 119 245 120 247 257 258 cell_2rw
* cell instance $1466 m0 *1 16.45,89.7
X$1466 117 118 119 250 120 249 257 258 cell_2rw
* cell instance $1467 r0 *1 16.45,89.7
X$1467 117 118 119 246 120 248 257 258 cell_2rw
* cell instance $1468 m0 *1 16.45,92.69
X$1468 117 118 119 253 120 256 257 258 cell_2rw
* cell instance $1469 r0 *1 16.45,92.69
X$1469 117 118 119 255 120 254 257 258 cell_2rw
* cell instance $1470 m0 *1 16.45,95.68
X$1470 117 118 119 251 120 252 257 258 cell_2rw
* cell instance $1471 r0 *1 17.625,44.85
X$1471 121 122 123 127 124 128 257 258 cell_2rw
* cell instance $1472 m0 *1 17.625,47.84
X$1472 121 122 123 126 124 125 257 258 cell_2rw
* cell instance $1473 m0 *1 17.625,50.83
X$1473 121 122 123 195 124 197 257 258 cell_2rw
* cell instance $1474 r0 *1 17.625,47.84
X$1474 121 122 123 199 124 201 257 258 cell_2rw
* cell instance $1475 r0 *1 17.625,50.83
X$1475 121 122 123 202 124 194 257 258 cell_2rw
* cell instance $1476 m0 *1 17.625,53.82
X$1476 121 122 123 198 124 193 257 258 cell_2rw
* cell instance $1477 m0 *1 17.625,56.81
X$1477 121 122 123 203 124 207 257 258 cell_2rw
* cell instance $1478 r0 *1 17.625,53.82
X$1478 121 122 123 196 124 200 257 258 cell_2rw
* cell instance $1479 m0 *1 17.625,59.8
X$1479 121 122 123 205 124 204 257 258 cell_2rw
* cell instance $1480 r0 *1 17.625,56.81
X$1480 121 122 123 206 124 208 257 258 cell_2rw
* cell instance $1481 m0 *1 17.625,62.79
X$1481 121 122 123 212 124 211 257 258 cell_2rw
* cell instance $1482 r0 *1 17.625,59.8
X$1482 121 122 123 214 124 213 257 258 cell_2rw
* cell instance $1483 m0 *1 17.625,65.78
X$1483 121 122 123 219 124 217 257 258 cell_2rw
* cell instance $1484 r0 *1 17.625,62.79
X$1484 121 122 123 210 124 209 257 258 cell_2rw
* cell instance $1485 r0 *1 17.625,65.78
X$1485 121 122 123 216 124 215 257 258 cell_2rw
* cell instance $1486 m0 *1 17.625,68.77
X$1486 121 122 123 218 124 220 257 258 cell_2rw
* cell instance $1487 m0 *1 17.625,71.76
X$1487 121 122 123 221 124 222 257 258 cell_2rw
* cell instance $1488 r0 *1 17.625,68.77
X$1488 121 122 123 224 124 223 257 258 cell_2rw
* cell instance $1489 r0 *1 17.625,71.76
X$1489 121 122 123 226 124 225 257 258 cell_2rw
* cell instance $1490 m0 *1 17.625,74.75
X$1490 121 122 123 231 124 232 257 258 cell_2rw
* cell instance $1491 r0 *1 17.625,74.75
X$1491 121 122 123 230 124 229 257 258 cell_2rw
* cell instance $1492 m0 *1 17.625,77.74
X$1492 121 122 123 227 124 228 257 258 cell_2rw
* cell instance $1493 r0 *1 17.625,77.74
X$1493 121 122 123 237 124 238 257 258 cell_2rw
* cell instance $1494 m0 *1 17.625,80.73
X$1494 121 122 123 233 124 236 257 258 cell_2rw
* cell instance $1495 r0 *1 17.625,80.73
X$1495 121 122 123 235 124 234 257 258 cell_2rw
* cell instance $1496 m0 *1 17.625,83.72
X$1496 121 122 123 240 124 242 257 258 cell_2rw
* cell instance $1497 r0 *1 17.625,83.72
X$1497 121 122 123 239 124 241 257 258 cell_2rw
* cell instance $1498 m0 *1 17.625,86.71
X$1498 121 122 123 244 124 243 257 258 cell_2rw
* cell instance $1499 r0 *1 17.625,86.71
X$1499 121 122 123 245 124 247 257 258 cell_2rw
* cell instance $1500 m0 *1 17.625,89.7
X$1500 121 122 123 250 124 249 257 258 cell_2rw
* cell instance $1501 m0 *1 17.625,92.69
X$1501 121 122 123 253 124 256 257 258 cell_2rw
* cell instance $1502 r0 *1 17.625,89.7
X$1502 121 122 123 246 124 248 257 258 cell_2rw
* cell instance $1503 m0 *1 17.625,95.68
X$1503 121 122 123 251 124 252 257 258 cell_2rw
* cell instance $1504 r0 *1 17.625,92.69
X$1504 121 122 123 255 124 254 257 258 cell_2rw
* cell instance $1505 m0 *1 18.8,47.84
X$1505 129 130 131 126 132 125 257 258 cell_2rw
* cell instance $1506 m0 *1 19.975,47.84
X$1506 133 134 135 126 136 125 257 258 cell_2rw
* cell instance $1507 m0 *1 21.15,47.84
X$1507 137 138 139 126 140 125 257 258 cell_2rw
* cell instance $1508 m0 *1 22.325,47.84
X$1508 141 142 143 126 144 125 257 258 cell_2rw
* cell instance $1509 m0 *1 23.5,47.84
X$1509 145 146 147 126 148 125 257 258 cell_2rw
* cell instance $1510 m0 *1 24.675,47.84
X$1510 149 150 151 126 152 125 257 258 cell_2rw
* cell instance $1511 m0 *1 25.85,47.84
X$1511 153 154 155 126 156 125 257 258 cell_2rw
* cell instance $1512 m0 *1 27.025,47.84
X$1512 157 158 159 126 160 125 257 258 cell_2rw
* cell instance $1513 m0 *1 28.2,47.84
X$1513 161 162 163 126 164 125 257 258 cell_2rw
* cell instance $1514 m0 *1 29.375,47.84
X$1514 165 166 167 126 168 125 257 258 cell_2rw
* cell instance $1515 m0 *1 30.55,47.84
X$1515 169 170 171 126 172 125 257 258 cell_2rw
* cell instance $1516 m0 *1 31.725,47.84
X$1516 173 174 175 126 176 125 257 258 cell_2rw
* cell instance $1517 m0 *1 32.9,47.84
X$1517 177 178 179 126 180 125 257 258 cell_2rw
* cell instance $1518 m0 *1 34.075,47.84
X$1518 181 182 183 126 184 125 257 258 cell_2rw
* cell instance $1519 m0 *1 35.25,47.84
X$1519 185 186 187 126 188 125 257 258 cell_2rw
* cell instance $1520 m0 *1 36.425,47.84
X$1520 189 190 191 126 192 125 257 258 cell_2rw
* cell instance $1521 r0 *1 18.8,44.85
X$1521 129 130 131 127 132 128 257 258 cell_2rw
* cell instance $1522 r0 *1 19.975,44.85
X$1522 133 134 135 127 136 128 257 258 cell_2rw
* cell instance $1523 r0 *1 21.15,44.85
X$1523 137 138 139 127 140 128 257 258 cell_2rw
* cell instance $1524 r0 *1 22.325,44.85
X$1524 141 142 143 127 144 128 257 258 cell_2rw
* cell instance $1525 r0 *1 23.5,44.85
X$1525 145 146 147 127 148 128 257 258 cell_2rw
* cell instance $1526 r0 *1 24.675,44.85
X$1526 149 150 151 127 152 128 257 258 cell_2rw
* cell instance $1527 r0 *1 25.85,44.85
X$1527 153 154 155 127 156 128 257 258 cell_2rw
* cell instance $1528 r0 *1 27.025,44.85
X$1528 157 158 159 127 160 128 257 258 cell_2rw
* cell instance $1529 r0 *1 28.2,44.85
X$1529 161 162 163 127 164 128 257 258 cell_2rw
* cell instance $1530 r0 *1 29.375,44.85
X$1530 165 166 167 127 168 128 257 258 cell_2rw
* cell instance $1531 r0 *1 30.55,44.85
X$1531 169 170 171 127 172 128 257 258 cell_2rw
* cell instance $1532 r0 *1 31.725,44.85
X$1532 173 174 175 127 176 128 257 258 cell_2rw
* cell instance $1533 r0 *1 32.9,44.85
X$1533 177 178 179 127 180 128 257 258 cell_2rw
* cell instance $1534 r0 *1 34.075,44.85
X$1534 181 182 183 127 184 128 257 258 cell_2rw
* cell instance $1535 r0 *1 35.25,44.85
X$1535 185 186 187 127 188 128 257 258 cell_2rw
* cell instance $1536 r0 *1 36.425,44.85
X$1536 189 190 191 127 192 128 257 258 cell_2rw
* cell instance $1537 r0 *1 18.8,47.84
X$1537 129 130 131 199 132 201 257 258 cell_2rw
* cell instance $1538 m0 *1 18.8,50.83
X$1538 129 130 131 195 132 197 257 258 cell_2rw
* cell instance $1539 r0 *1 18.8,50.83
X$1539 129 130 131 202 132 194 257 258 cell_2rw
* cell instance $1540 m0 *1 18.8,53.82
X$1540 129 130 131 198 132 193 257 258 cell_2rw
* cell instance $1541 r0 *1 18.8,53.82
X$1541 129 130 131 196 132 200 257 258 cell_2rw
* cell instance $1542 m0 *1 18.8,56.81
X$1542 129 130 131 203 132 207 257 258 cell_2rw
* cell instance $1543 r0 *1 18.8,56.81
X$1543 129 130 131 206 132 208 257 258 cell_2rw
* cell instance $1544 m0 *1 18.8,59.8
X$1544 129 130 131 205 132 204 257 258 cell_2rw
* cell instance $1545 r0 *1 18.8,59.8
X$1545 129 130 131 214 132 213 257 258 cell_2rw
* cell instance $1546 m0 *1 18.8,62.79
X$1546 129 130 131 212 132 211 257 258 cell_2rw
* cell instance $1547 r0 *1 18.8,62.79
X$1547 129 130 131 210 132 209 257 258 cell_2rw
* cell instance $1548 m0 *1 18.8,65.78
X$1548 129 130 131 219 132 217 257 258 cell_2rw
* cell instance $1549 r0 *1 18.8,65.78
X$1549 129 130 131 216 132 215 257 258 cell_2rw
* cell instance $1550 m0 *1 18.8,68.77
X$1550 129 130 131 218 132 220 257 258 cell_2rw
* cell instance $1551 m0 *1 18.8,71.76
X$1551 129 130 131 221 132 222 257 258 cell_2rw
* cell instance $1552 r0 *1 18.8,68.77
X$1552 129 130 131 224 132 223 257 258 cell_2rw
* cell instance $1553 m0 *1 18.8,74.75
X$1553 129 130 131 231 132 232 257 258 cell_2rw
* cell instance $1554 r0 *1 18.8,71.76
X$1554 129 130 131 226 132 225 257 258 cell_2rw
* cell instance $1555 m0 *1 18.8,77.74
X$1555 129 130 131 227 132 228 257 258 cell_2rw
* cell instance $1556 r0 *1 18.8,74.75
X$1556 129 130 131 230 132 229 257 258 cell_2rw
* cell instance $1557 r0 *1 18.8,77.74
X$1557 129 130 131 237 132 238 257 258 cell_2rw
* cell instance $1558 m0 *1 18.8,80.73
X$1558 129 130 131 233 132 236 257 258 cell_2rw
* cell instance $1559 r0 *1 18.8,80.73
X$1559 129 130 131 235 132 234 257 258 cell_2rw
* cell instance $1560 m0 *1 18.8,83.72
X$1560 129 130 131 240 132 242 257 258 cell_2rw
* cell instance $1561 r0 *1 18.8,83.72
X$1561 129 130 131 239 132 241 257 258 cell_2rw
* cell instance $1562 m0 *1 18.8,86.71
X$1562 129 130 131 244 132 243 257 258 cell_2rw
* cell instance $1563 r0 *1 18.8,86.71
X$1563 129 130 131 245 132 247 257 258 cell_2rw
* cell instance $1564 m0 *1 18.8,89.7
X$1564 129 130 131 250 132 249 257 258 cell_2rw
* cell instance $1565 r0 *1 18.8,89.7
X$1565 129 130 131 246 132 248 257 258 cell_2rw
* cell instance $1566 m0 *1 18.8,92.69
X$1566 129 130 131 253 132 256 257 258 cell_2rw
* cell instance $1567 r0 *1 18.8,92.69
X$1567 129 130 131 255 132 254 257 258 cell_2rw
* cell instance $1568 m0 *1 18.8,95.68
X$1568 129 130 131 251 132 252 257 258 cell_2rw
* cell instance $1569 r0 *1 19.975,47.84
X$1569 133 134 135 199 136 201 257 258 cell_2rw
* cell instance $1570 m0 *1 19.975,50.83
X$1570 133 134 135 195 136 197 257 258 cell_2rw
* cell instance $1571 r0 *1 19.975,50.83
X$1571 133 134 135 202 136 194 257 258 cell_2rw
* cell instance $1572 m0 *1 19.975,53.82
X$1572 133 134 135 198 136 193 257 258 cell_2rw
* cell instance $1573 m0 *1 19.975,56.81
X$1573 133 134 135 203 136 207 257 258 cell_2rw
* cell instance $1574 r0 *1 19.975,53.82
X$1574 133 134 135 196 136 200 257 258 cell_2rw
* cell instance $1575 r0 *1 19.975,56.81
X$1575 133 134 135 206 136 208 257 258 cell_2rw
* cell instance $1576 m0 *1 19.975,59.8
X$1576 133 134 135 205 136 204 257 258 cell_2rw
* cell instance $1577 r0 *1 19.975,59.8
X$1577 133 134 135 214 136 213 257 258 cell_2rw
* cell instance $1578 m0 *1 19.975,62.79
X$1578 133 134 135 212 136 211 257 258 cell_2rw
* cell instance $1579 r0 *1 19.975,62.79
X$1579 133 134 135 210 136 209 257 258 cell_2rw
* cell instance $1580 m0 *1 19.975,65.78
X$1580 133 134 135 219 136 217 257 258 cell_2rw
* cell instance $1581 r0 *1 19.975,65.78
X$1581 133 134 135 216 136 215 257 258 cell_2rw
* cell instance $1582 m0 *1 19.975,68.77
X$1582 133 134 135 218 136 220 257 258 cell_2rw
* cell instance $1583 r0 *1 19.975,68.77
X$1583 133 134 135 224 136 223 257 258 cell_2rw
* cell instance $1584 m0 *1 19.975,71.76
X$1584 133 134 135 221 136 222 257 258 cell_2rw
* cell instance $1585 r0 *1 19.975,71.76
X$1585 133 134 135 226 136 225 257 258 cell_2rw
* cell instance $1586 m0 *1 19.975,74.75
X$1586 133 134 135 231 136 232 257 258 cell_2rw
* cell instance $1587 r0 *1 19.975,74.75
X$1587 133 134 135 230 136 229 257 258 cell_2rw
* cell instance $1588 m0 *1 19.975,77.74
X$1588 133 134 135 227 136 228 257 258 cell_2rw
* cell instance $1589 m0 *1 19.975,80.73
X$1589 133 134 135 233 136 236 257 258 cell_2rw
* cell instance $1590 r0 *1 19.975,77.74
X$1590 133 134 135 237 136 238 257 258 cell_2rw
* cell instance $1591 r0 *1 19.975,80.73
X$1591 133 134 135 235 136 234 257 258 cell_2rw
* cell instance $1592 m0 *1 19.975,83.72
X$1592 133 134 135 240 136 242 257 258 cell_2rw
* cell instance $1593 r0 *1 19.975,83.72
X$1593 133 134 135 239 136 241 257 258 cell_2rw
* cell instance $1594 m0 *1 19.975,86.71
X$1594 133 134 135 244 136 243 257 258 cell_2rw
* cell instance $1595 r0 *1 19.975,86.71
X$1595 133 134 135 245 136 247 257 258 cell_2rw
* cell instance $1596 m0 *1 19.975,89.7
X$1596 133 134 135 250 136 249 257 258 cell_2rw
* cell instance $1597 r0 *1 19.975,89.7
X$1597 133 134 135 246 136 248 257 258 cell_2rw
* cell instance $1598 m0 *1 19.975,92.69
X$1598 133 134 135 253 136 256 257 258 cell_2rw
* cell instance $1599 r0 *1 19.975,92.69
X$1599 133 134 135 255 136 254 257 258 cell_2rw
* cell instance $1600 m0 *1 19.975,95.68
X$1600 133 134 135 251 136 252 257 258 cell_2rw
* cell instance $1601 r0 *1 21.15,47.84
X$1601 137 138 139 199 140 201 257 258 cell_2rw
* cell instance $1602 m0 *1 21.15,50.83
X$1602 137 138 139 195 140 197 257 258 cell_2rw
* cell instance $1603 r0 *1 21.15,50.83
X$1603 137 138 139 202 140 194 257 258 cell_2rw
* cell instance $1604 m0 *1 21.15,53.82
X$1604 137 138 139 198 140 193 257 258 cell_2rw
* cell instance $1605 r0 *1 21.15,53.82
X$1605 137 138 139 196 140 200 257 258 cell_2rw
* cell instance $1606 m0 *1 21.15,56.81
X$1606 137 138 139 203 140 207 257 258 cell_2rw
* cell instance $1607 r0 *1 21.15,56.81
X$1607 137 138 139 206 140 208 257 258 cell_2rw
* cell instance $1608 m0 *1 21.15,59.8
X$1608 137 138 139 205 140 204 257 258 cell_2rw
* cell instance $1609 r0 *1 21.15,59.8
X$1609 137 138 139 214 140 213 257 258 cell_2rw
* cell instance $1610 m0 *1 21.15,62.79
X$1610 137 138 139 212 140 211 257 258 cell_2rw
* cell instance $1611 r0 *1 21.15,62.79
X$1611 137 138 139 210 140 209 257 258 cell_2rw
* cell instance $1612 m0 *1 21.15,65.78
X$1612 137 138 139 219 140 217 257 258 cell_2rw
* cell instance $1613 r0 *1 21.15,65.78
X$1613 137 138 139 216 140 215 257 258 cell_2rw
* cell instance $1614 m0 *1 21.15,68.77
X$1614 137 138 139 218 140 220 257 258 cell_2rw
* cell instance $1615 r0 *1 21.15,68.77
X$1615 137 138 139 224 140 223 257 258 cell_2rw
* cell instance $1616 m0 *1 21.15,71.76
X$1616 137 138 139 221 140 222 257 258 cell_2rw
* cell instance $1617 r0 *1 21.15,71.76
X$1617 137 138 139 226 140 225 257 258 cell_2rw
* cell instance $1618 m0 *1 21.15,74.75
X$1618 137 138 139 231 140 232 257 258 cell_2rw
* cell instance $1619 r0 *1 21.15,74.75
X$1619 137 138 139 230 140 229 257 258 cell_2rw
* cell instance $1620 m0 *1 21.15,77.74
X$1620 137 138 139 227 140 228 257 258 cell_2rw
* cell instance $1621 r0 *1 21.15,77.74
X$1621 137 138 139 237 140 238 257 258 cell_2rw
* cell instance $1622 m0 *1 21.15,80.73
X$1622 137 138 139 233 140 236 257 258 cell_2rw
* cell instance $1623 r0 *1 21.15,80.73
X$1623 137 138 139 235 140 234 257 258 cell_2rw
* cell instance $1624 m0 *1 21.15,83.72
X$1624 137 138 139 240 140 242 257 258 cell_2rw
* cell instance $1625 r0 *1 21.15,83.72
X$1625 137 138 139 239 140 241 257 258 cell_2rw
* cell instance $1626 m0 *1 21.15,86.71
X$1626 137 138 139 244 140 243 257 258 cell_2rw
* cell instance $1627 r0 *1 21.15,86.71
X$1627 137 138 139 245 140 247 257 258 cell_2rw
* cell instance $1628 m0 *1 21.15,89.7
X$1628 137 138 139 250 140 249 257 258 cell_2rw
* cell instance $1629 r0 *1 21.15,89.7
X$1629 137 138 139 246 140 248 257 258 cell_2rw
* cell instance $1630 m0 *1 21.15,92.69
X$1630 137 138 139 253 140 256 257 258 cell_2rw
* cell instance $1631 r0 *1 21.15,92.69
X$1631 137 138 139 255 140 254 257 258 cell_2rw
* cell instance $1632 m0 *1 21.15,95.68
X$1632 137 138 139 251 140 252 257 258 cell_2rw
* cell instance $1633 r0 *1 22.325,47.84
X$1633 141 142 143 199 144 201 257 258 cell_2rw
* cell instance $1634 m0 *1 22.325,50.83
X$1634 141 142 143 195 144 197 257 258 cell_2rw
* cell instance $1635 r0 *1 22.325,50.83
X$1635 141 142 143 202 144 194 257 258 cell_2rw
* cell instance $1636 m0 *1 22.325,53.82
X$1636 141 142 143 198 144 193 257 258 cell_2rw
* cell instance $1637 m0 *1 22.325,56.81
X$1637 141 142 143 203 144 207 257 258 cell_2rw
* cell instance $1638 r0 *1 22.325,53.82
X$1638 141 142 143 196 144 200 257 258 cell_2rw
* cell instance $1639 r0 *1 22.325,56.81
X$1639 141 142 143 206 144 208 257 258 cell_2rw
* cell instance $1640 m0 *1 22.325,59.8
X$1640 141 142 143 205 144 204 257 258 cell_2rw
* cell instance $1641 r0 *1 22.325,59.8
X$1641 141 142 143 214 144 213 257 258 cell_2rw
* cell instance $1642 m0 *1 22.325,62.79
X$1642 141 142 143 212 144 211 257 258 cell_2rw
* cell instance $1643 r0 *1 22.325,62.79
X$1643 141 142 143 210 144 209 257 258 cell_2rw
* cell instance $1644 m0 *1 22.325,65.78
X$1644 141 142 143 219 144 217 257 258 cell_2rw
* cell instance $1645 r0 *1 22.325,65.78
X$1645 141 142 143 216 144 215 257 258 cell_2rw
* cell instance $1646 m0 *1 22.325,68.77
X$1646 141 142 143 218 144 220 257 258 cell_2rw
* cell instance $1647 r0 *1 22.325,68.77
X$1647 141 142 143 224 144 223 257 258 cell_2rw
* cell instance $1648 m0 *1 22.325,71.76
X$1648 141 142 143 221 144 222 257 258 cell_2rw
* cell instance $1649 r0 *1 22.325,71.76
X$1649 141 142 143 226 144 225 257 258 cell_2rw
* cell instance $1650 m0 *1 22.325,74.75
X$1650 141 142 143 231 144 232 257 258 cell_2rw
* cell instance $1651 r0 *1 22.325,74.75
X$1651 141 142 143 230 144 229 257 258 cell_2rw
* cell instance $1652 m0 *1 22.325,77.74
X$1652 141 142 143 227 144 228 257 258 cell_2rw
* cell instance $1653 r0 *1 22.325,77.74
X$1653 141 142 143 237 144 238 257 258 cell_2rw
* cell instance $1654 m0 *1 22.325,80.73
X$1654 141 142 143 233 144 236 257 258 cell_2rw
* cell instance $1655 r0 *1 22.325,80.73
X$1655 141 142 143 235 144 234 257 258 cell_2rw
* cell instance $1656 m0 *1 22.325,83.72
X$1656 141 142 143 240 144 242 257 258 cell_2rw
* cell instance $1657 r0 *1 22.325,83.72
X$1657 141 142 143 239 144 241 257 258 cell_2rw
* cell instance $1658 m0 *1 22.325,86.71
X$1658 141 142 143 244 144 243 257 258 cell_2rw
* cell instance $1659 m0 *1 22.325,89.7
X$1659 141 142 143 250 144 249 257 258 cell_2rw
* cell instance $1660 r0 *1 22.325,86.71
X$1660 141 142 143 245 144 247 257 258 cell_2rw
* cell instance $1661 m0 *1 22.325,92.69
X$1661 141 142 143 253 144 256 257 258 cell_2rw
* cell instance $1662 r0 *1 22.325,89.7
X$1662 141 142 143 246 144 248 257 258 cell_2rw
* cell instance $1663 r0 *1 22.325,92.69
X$1663 141 142 143 255 144 254 257 258 cell_2rw
* cell instance $1664 m0 *1 22.325,95.68
X$1664 141 142 143 251 144 252 257 258 cell_2rw
* cell instance $1665 r0 *1 23.5,47.84
X$1665 145 146 147 199 148 201 257 258 cell_2rw
* cell instance $1666 m0 *1 23.5,50.83
X$1666 145 146 147 195 148 197 257 258 cell_2rw
* cell instance $1667 r0 *1 23.5,50.83
X$1667 145 146 147 202 148 194 257 258 cell_2rw
* cell instance $1668 m0 *1 23.5,53.82
X$1668 145 146 147 198 148 193 257 258 cell_2rw
* cell instance $1669 r0 *1 23.5,53.82
X$1669 145 146 147 196 148 200 257 258 cell_2rw
* cell instance $1670 m0 *1 23.5,56.81
X$1670 145 146 147 203 148 207 257 258 cell_2rw
* cell instance $1671 r0 *1 23.5,56.81
X$1671 145 146 147 206 148 208 257 258 cell_2rw
* cell instance $1672 m0 *1 23.5,59.8
X$1672 145 146 147 205 148 204 257 258 cell_2rw
* cell instance $1673 r0 *1 23.5,59.8
X$1673 145 146 147 214 148 213 257 258 cell_2rw
* cell instance $1674 m0 *1 23.5,62.79
X$1674 145 146 147 212 148 211 257 258 cell_2rw
* cell instance $1675 r0 *1 23.5,62.79
X$1675 145 146 147 210 148 209 257 258 cell_2rw
* cell instance $1676 m0 *1 23.5,65.78
X$1676 145 146 147 219 148 217 257 258 cell_2rw
* cell instance $1677 r0 *1 23.5,65.78
X$1677 145 146 147 216 148 215 257 258 cell_2rw
* cell instance $1678 m0 *1 23.5,68.77
X$1678 145 146 147 218 148 220 257 258 cell_2rw
* cell instance $1679 m0 *1 23.5,71.76
X$1679 145 146 147 221 148 222 257 258 cell_2rw
* cell instance $1680 r0 *1 23.5,68.77
X$1680 145 146 147 224 148 223 257 258 cell_2rw
* cell instance $1681 r0 *1 23.5,71.76
X$1681 145 146 147 226 148 225 257 258 cell_2rw
* cell instance $1682 m0 *1 23.5,74.75
X$1682 145 146 147 231 148 232 257 258 cell_2rw
* cell instance $1683 r0 *1 23.5,74.75
X$1683 145 146 147 230 148 229 257 258 cell_2rw
* cell instance $1684 m0 *1 23.5,77.74
X$1684 145 146 147 227 148 228 257 258 cell_2rw
* cell instance $1685 r0 *1 23.5,77.74
X$1685 145 146 147 237 148 238 257 258 cell_2rw
* cell instance $1686 m0 *1 23.5,80.73
X$1686 145 146 147 233 148 236 257 258 cell_2rw
* cell instance $1687 m0 *1 23.5,83.72
X$1687 145 146 147 240 148 242 257 258 cell_2rw
* cell instance $1688 r0 *1 23.5,80.73
X$1688 145 146 147 235 148 234 257 258 cell_2rw
* cell instance $1689 r0 *1 23.5,83.72
X$1689 145 146 147 239 148 241 257 258 cell_2rw
* cell instance $1690 m0 *1 23.5,86.71
X$1690 145 146 147 244 148 243 257 258 cell_2rw
* cell instance $1691 r0 *1 23.5,86.71
X$1691 145 146 147 245 148 247 257 258 cell_2rw
* cell instance $1692 m0 *1 23.5,89.7
X$1692 145 146 147 250 148 249 257 258 cell_2rw
* cell instance $1693 r0 *1 23.5,89.7
X$1693 145 146 147 246 148 248 257 258 cell_2rw
* cell instance $1694 m0 *1 23.5,92.69
X$1694 145 146 147 253 148 256 257 258 cell_2rw
* cell instance $1695 m0 *1 23.5,95.68
X$1695 145 146 147 251 148 252 257 258 cell_2rw
* cell instance $1696 r0 *1 23.5,92.69
X$1696 145 146 147 255 148 254 257 258 cell_2rw
* cell instance $1697 r0 *1 24.675,47.84
X$1697 149 150 151 199 152 201 257 258 cell_2rw
* cell instance $1698 m0 *1 24.675,50.83
X$1698 149 150 151 195 152 197 257 258 cell_2rw
* cell instance $1699 r0 *1 24.675,50.83
X$1699 149 150 151 202 152 194 257 258 cell_2rw
* cell instance $1700 m0 *1 24.675,53.82
X$1700 149 150 151 198 152 193 257 258 cell_2rw
* cell instance $1701 r0 *1 24.675,53.82
X$1701 149 150 151 196 152 200 257 258 cell_2rw
* cell instance $1702 m0 *1 24.675,56.81
X$1702 149 150 151 203 152 207 257 258 cell_2rw
* cell instance $1703 r0 *1 24.675,56.81
X$1703 149 150 151 206 152 208 257 258 cell_2rw
* cell instance $1704 m0 *1 24.675,59.8
X$1704 149 150 151 205 152 204 257 258 cell_2rw
* cell instance $1705 r0 *1 24.675,59.8
X$1705 149 150 151 214 152 213 257 258 cell_2rw
* cell instance $1706 m0 *1 24.675,62.79
X$1706 149 150 151 212 152 211 257 258 cell_2rw
* cell instance $1707 r0 *1 24.675,62.79
X$1707 149 150 151 210 152 209 257 258 cell_2rw
* cell instance $1708 m0 *1 24.675,65.78
X$1708 149 150 151 219 152 217 257 258 cell_2rw
* cell instance $1709 r0 *1 24.675,65.78
X$1709 149 150 151 216 152 215 257 258 cell_2rw
* cell instance $1710 m0 *1 24.675,68.77
X$1710 149 150 151 218 152 220 257 258 cell_2rw
* cell instance $1711 r0 *1 24.675,68.77
X$1711 149 150 151 224 152 223 257 258 cell_2rw
* cell instance $1712 m0 *1 24.675,71.76
X$1712 149 150 151 221 152 222 257 258 cell_2rw
* cell instance $1713 m0 *1 24.675,74.75
X$1713 149 150 151 231 152 232 257 258 cell_2rw
* cell instance $1714 r0 *1 24.675,71.76
X$1714 149 150 151 226 152 225 257 258 cell_2rw
* cell instance $1715 r0 *1 24.675,74.75
X$1715 149 150 151 230 152 229 257 258 cell_2rw
* cell instance $1716 m0 *1 24.675,77.74
X$1716 149 150 151 227 152 228 257 258 cell_2rw
* cell instance $1717 r0 *1 24.675,77.74
X$1717 149 150 151 237 152 238 257 258 cell_2rw
* cell instance $1718 m0 *1 24.675,80.73
X$1718 149 150 151 233 152 236 257 258 cell_2rw
* cell instance $1719 r0 *1 24.675,80.73
X$1719 149 150 151 235 152 234 257 258 cell_2rw
* cell instance $1720 m0 *1 24.675,83.72
X$1720 149 150 151 240 152 242 257 258 cell_2rw
* cell instance $1721 r0 *1 24.675,83.72
X$1721 149 150 151 239 152 241 257 258 cell_2rw
* cell instance $1722 m0 *1 24.675,86.71
X$1722 149 150 151 244 152 243 257 258 cell_2rw
* cell instance $1723 r0 *1 24.675,86.71
X$1723 149 150 151 245 152 247 257 258 cell_2rw
* cell instance $1724 m0 *1 24.675,89.7
X$1724 149 150 151 250 152 249 257 258 cell_2rw
* cell instance $1725 r0 *1 24.675,89.7
X$1725 149 150 151 246 152 248 257 258 cell_2rw
* cell instance $1726 m0 *1 24.675,92.69
X$1726 149 150 151 253 152 256 257 258 cell_2rw
* cell instance $1727 m0 *1 24.675,95.68
X$1727 149 150 151 251 152 252 257 258 cell_2rw
* cell instance $1728 r0 *1 24.675,92.69
X$1728 149 150 151 255 152 254 257 258 cell_2rw
* cell instance $1729 r0 *1 25.85,47.84
X$1729 153 154 155 199 156 201 257 258 cell_2rw
* cell instance $1730 m0 *1 25.85,50.83
X$1730 153 154 155 195 156 197 257 258 cell_2rw
* cell instance $1731 r0 *1 25.85,50.83
X$1731 153 154 155 202 156 194 257 258 cell_2rw
* cell instance $1732 m0 *1 25.85,53.82
X$1732 153 154 155 198 156 193 257 258 cell_2rw
* cell instance $1733 r0 *1 25.85,53.82
X$1733 153 154 155 196 156 200 257 258 cell_2rw
* cell instance $1734 m0 *1 25.85,56.81
X$1734 153 154 155 203 156 207 257 258 cell_2rw
* cell instance $1735 r0 *1 25.85,56.81
X$1735 153 154 155 206 156 208 257 258 cell_2rw
* cell instance $1736 m0 *1 25.85,59.8
X$1736 153 154 155 205 156 204 257 258 cell_2rw
* cell instance $1737 r0 *1 25.85,59.8
X$1737 153 154 155 214 156 213 257 258 cell_2rw
* cell instance $1738 m0 *1 25.85,62.79
X$1738 153 154 155 212 156 211 257 258 cell_2rw
* cell instance $1739 m0 *1 25.85,65.78
X$1739 153 154 155 219 156 217 257 258 cell_2rw
* cell instance $1740 r0 *1 25.85,62.79
X$1740 153 154 155 210 156 209 257 258 cell_2rw
* cell instance $1741 r0 *1 25.85,65.78
X$1741 153 154 155 216 156 215 257 258 cell_2rw
* cell instance $1742 m0 *1 25.85,68.77
X$1742 153 154 155 218 156 220 257 258 cell_2rw
* cell instance $1743 m0 *1 25.85,71.76
X$1743 153 154 155 221 156 222 257 258 cell_2rw
* cell instance $1744 r0 *1 25.85,68.77
X$1744 153 154 155 224 156 223 257 258 cell_2rw
* cell instance $1745 r0 *1 25.85,71.76
X$1745 153 154 155 226 156 225 257 258 cell_2rw
* cell instance $1746 m0 *1 25.85,74.75
X$1746 153 154 155 231 156 232 257 258 cell_2rw
* cell instance $1747 r0 *1 25.85,74.75
X$1747 153 154 155 230 156 229 257 258 cell_2rw
* cell instance $1748 m0 *1 25.85,77.74
X$1748 153 154 155 227 156 228 257 258 cell_2rw
* cell instance $1749 r0 *1 25.85,77.74
X$1749 153 154 155 237 156 238 257 258 cell_2rw
* cell instance $1750 m0 *1 25.85,80.73
X$1750 153 154 155 233 156 236 257 258 cell_2rw
* cell instance $1751 r0 *1 25.85,80.73
X$1751 153 154 155 235 156 234 257 258 cell_2rw
* cell instance $1752 m0 *1 25.85,83.72
X$1752 153 154 155 240 156 242 257 258 cell_2rw
* cell instance $1753 r0 *1 25.85,83.72
X$1753 153 154 155 239 156 241 257 258 cell_2rw
* cell instance $1754 m0 *1 25.85,86.71
X$1754 153 154 155 244 156 243 257 258 cell_2rw
* cell instance $1755 r0 *1 25.85,86.71
X$1755 153 154 155 245 156 247 257 258 cell_2rw
* cell instance $1756 m0 *1 25.85,89.7
X$1756 153 154 155 250 156 249 257 258 cell_2rw
* cell instance $1757 r0 *1 25.85,89.7
X$1757 153 154 155 246 156 248 257 258 cell_2rw
* cell instance $1758 m0 *1 25.85,92.69
X$1758 153 154 155 253 156 256 257 258 cell_2rw
* cell instance $1759 m0 *1 25.85,95.68
X$1759 153 154 155 251 156 252 257 258 cell_2rw
* cell instance $1760 r0 *1 25.85,92.69
X$1760 153 154 155 255 156 254 257 258 cell_2rw
* cell instance $1761 r0 *1 27.025,47.84
X$1761 157 158 159 199 160 201 257 258 cell_2rw
* cell instance $1762 m0 *1 27.025,50.83
X$1762 157 158 159 195 160 197 257 258 cell_2rw
* cell instance $1763 m0 *1 27.025,53.82
X$1763 157 158 159 198 160 193 257 258 cell_2rw
* cell instance $1764 r0 *1 27.025,50.83
X$1764 157 158 159 202 160 194 257 258 cell_2rw
* cell instance $1765 m0 *1 27.025,56.81
X$1765 157 158 159 203 160 207 257 258 cell_2rw
* cell instance $1766 r0 *1 27.025,53.82
X$1766 157 158 159 196 160 200 257 258 cell_2rw
* cell instance $1767 r0 *1 27.025,56.81
X$1767 157 158 159 206 160 208 257 258 cell_2rw
* cell instance $1768 m0 *1 27.025,59.8
X$1768 157 158 159 205 160 204 257 258 cell_2rw
* cell instance $1769 r0 *1 27.025,59.8
X$1769 157 158 159 214 160 213 257 258 cell_2rw
* cell instance $1770 m0 *1 27.025,62.79
X$1770 157 158 159 212 160 211 257 258 cell_2rw
* cell instance $1771 m0 *1 27.025,65.78
X$1771 157 158 159 219 160 217 257 258 cell_2rw
* cell instance $1772 r0 *1 27.025,62.79
X$1772 157 158 159 210 160 209 257 258 cell_2rw
* cell instance $1773 r0 *1 27.025,65.78
X$1773 157 158 159 216 160 215 257 258 cell_2rw
* cell instance $1774 m0 *1 27.025,68.77
X$1774 157 158 159 218 160 220 257 258 cell_2rw
* cell instance $1775 r0 *1 27.025,68.77
X$1775 157 158 159 224 160 223 257 258 cell_2rw
* cell instance $1776 m0 *1 27.025,71.76
X$1776 157 158 159 221 160 222 257 258 cell_2rw
* cell instance $1777 r0 *1 27.025,71.76
X$1777 157 158 159 226 160 225 257 258 cell_2rw
* cell instance $1778 m0 *1 27.025,74.75
X$1778 157 158 159 231 160 232 257 258 cell_2rw
* cell instance $1779 r0 *1 27.025,74.75
X$1779 157 158 159 230 160 229 257 258 cell_2rw
* cell instance $1780 m0 *1 27.025,77.74
X$1780 157 158 159 227 160 228 257 258 cell_2rw
* cell instance $1781 m0 *1 27.025,80.73
X$1781 157 158 159 233 160 236 257 258 cell_2rw
* cell instance $1782 r0 *1 27.025,77.74
X$1782 157 158 159 237 160 238 257 258 cell_2rw
* cell instance $1783 r0 *1 27.025,80.73
X$1783 157 158 159 235 160 234 257 258 cell_2rw
* cell instance $1784 m0 *1 27.025,83.72
X$1784 157 158 159 240 160 242 257 258 cell_2rw
* cell instance $1785 r0 *1 27.025,83.72
X$1785 157 158 159 239 160 241 257 258 cell_2rw
* cell instance $1786 m0 *1 27.025,86.71
X$1786 157 158 159 244 160 243 257 258 cell_2rw
* cell instance $1787 r0 *1 27.025,86.71
X$1787 157 158 159 245 160 247 257 258 cell_2rw
* cell instance $1788 m0 *1 27.025,89.7
X$1788 157 158 159 250 160 249 257 258 cell_2rw
* cell instance $1789 r0 *1 27.025,89.7
X$1789 157 158 159 246 160 248 257 258 cell_2rw
* cell instance $1790 m0 *1 27.025,92.69
X$1790 157 158 159 253 160 256 257 258 cell_2rw
* cell instance $1791 r0 *1 27.025,92.69
X$1791 157 158 159 255 160 254 257 258 cell_2rw
* cell instance $1792 m0 *1 27.025,95.68
X$1792 157 158 159 251 160 252 257 258 cell_2rw
* cell instance $1793 r0 *1 28.2,47.84
X$1793 161 162 163 199 164 201 257 258 cell_2rw
* cell instance $1794 m0 *1 28.2,50.83
X$1794 161 162 163 195 164 197 257 258 cell_2rw
* cell instance $1795 r0 *1 28.2,50.83
X$1795 161 162 163 202 164 194 257 258 cell_2rw
* cell instance $1796 m0 *1 28.2,53.82
X$1796 161 162 163 198 164 193 257 258 cell_2rw
* cell instance $1797 r0 *1 28.2,53.82
X$1797 161 162 163 196 164 200 257 258 cell_2rw
* cell instance $1798 m0 *1 28.2,56.81
X$1798 161 162 163 203 164 207 257 258 cell_2rw
* cell instance $1799 r0 *1 28.2,56.81
X$1799 161 162 163 206 164 208 257 258 cell_2rw
* cell instance $1800 m0 *1 28.2,59.8
X$1800 161 162 163 205 164 204 257 258 cell_2rw
* cell instance $1801 r0 *1 28.2,59.8
X$1801 161 162 163 214 164 213 257 258 cell_2rw
* cell instance $1802 m0 *1 28.2,62.79
X$1802 161 162 163 212 164 211 257 258 cell_2rw
* cell instance $1803 m0 *1 28.2,65.78
X$1803 161 162 163 219 164 217 257 258 cell_2rw
* cell instance $1804 r0 *1 28.2,62.79
X$1804 161 162 163 210 164 209 257 258 cell_2rw
* cell instance $1805 m0 *1 28.2,68.77
X$1805 161 162 163 218 164 220 257 258 cell_2rw
* cell instance $1806 r0 *1 28.2,65.78
X$1806 161 162 163 216 164 215 257 258 cell_2rw
* cell instance $1807 r0 *1 28.2,68.77
X$1807 161 162 163 224 164 223 257 258 cell_2rw
* cell instance $1808 m0 *1 28.2,71.76
X$1808 161 162 163 221 164 222 257 258 cell_2rw
* cell instance $1809 r0 *1 28.2,71.76
X$1809 161 162 163 226 164 225 257 258 cell_2rw
* cell instance $1810 m0 *1 28.2,74.75
X$1810 161 162 163 231 164 232 257 258 cell_2rw
* cell instance $1811 r0 *1 28.2,74.75
X$1811 161 162 163 230 164 229 257 258 cell_2rw
* cell instance $1812 m0 *1 28.2,77.74
X$1812 161 162 163 227 164 228 257 258 cell_2rw
* cell instance $1813 r0 *1 28.2,77.74
X$1813 161 162 163 237 164 238 257 258 cell_2rw
* cell instance $1814 m0 *1 28.2,80.73
X$1814 161 162 163 233 164 236 257 258 cell_2rw
* cell instance $1815 r0 *1 28.2,80.73
X$1815 161 162 163 235 164 234 257 258 cell_2rw
* cell instance $1816 m0 *1 28.2,83.72
X$1816 161 162 163 240 164 242 257 258 cell_2rw
* cell instance $1817 m0 *1 28.2,86.71
X$1817 161 162 163 244 164 243 257 258 cell_2rw
* cell instance $1818 r0 *1 28.2,83.72
X$1818 161 162 163 239 164 241 257 258 cell_2rw
* cell instance $1819 r0 *1 28.2,86.71
X$1819 161 162 163 245 164 247 257 258 cell_2rw
* cell instance $1820 m0 *1 28.2,89.7
X$1820 161 162 163 250 164 249 257 258 cell_2rw
* cell instance $1821 r0 *1 28.2,89.7
X$1821 161 162 163 246 164 248 257 258 cell_2rw
* cell instance $1822 m0 *1 28.2,92.69
X$1822 161 162 163 253 164 256 257 258 cell_2rw
* cell instance $1823 r0 *1 28.2,92.69
X$1823 161 162 163 255 164 254 257 258 cell_2rw
* cell instance $1824 m0 *1 28.2,95.68
X$1824 161 162 163 251 164 252 257 258 cell_2rw
* cell instance $1825 r0 *1 29.375,47.84
X$1825 165 166 167 199 168 201 257 258 cell_2rw
* cell instance $1826 m0 *1 29.375,50.83
X$1826 165 166 167 195 168 197 257 258 cell_2rw
* cell instance $1827 r0 *1 29.375,50.83
X$1827 165 166 167 202 168 194 257 258 cell_2rw
* cell instance $1828 m0 *1 29.375,53.82
X$1828 165 166 167 198 168 193 257 258 cell_2rw
* cell instance $1829 r0 *1 29.375,53.82
X$1829 165 166 167 196 168 200 257 258 cell_2rw
* cell instance $1830 m0 *1 29.375,56.81
X$1830 165 166 167 203 168 207 257 258 cell_2rw
* cell instance $1831 r0 *1 29.375,56.81
X$1831 165 166 167 206 168 208 257 258 cell_2rw
* cell instance $1832 m0 *1 29.375,59.8
X$1832 165 166 167 205 168 204 257 258 cell_2rw
* cell instance $1833 r0 *1 29.375,59.8
X$1833 165 166 167 214 168 213 257 258 cell_2rw
* cell instance $1834 m0 *1 29.375,62.79
X$1834 165 166 167 212 168 211 257 258 cell_2rw
* cell instance $1835 r0 *1 29.375,62.79
X$1835 165 166 167 210 168 209 257 258 cell_2rw
* cell instance $1836 m0 *1 29.375,65.78
X$1836 165 166 167 219 168 217 257 258 cell_2rw
* cell instance $1837 r0 *1 29.375,65.78
X$1837 165 166 167 216 168 215 257 258 cell_2rw
* cell instance $1838 m0 *1 29.375,68.77
X$1838 165 166 167 218 168 220 257 258 cell_2rw
* cell instance $1839 m0 *1 29.375,71.76
X$1839 165 166 167 221 168 222 257 258 cell_2rw
* cell instance $1840 r0 *1 29.375,68.77
X$1840 165 166 167 224 168 223 257 258 cell_2rw
* cell instance $1841 r0 *1 29.375,71.76
X$1841 165 166 167 226 168 225 257 258 cell_2rw
* cell instance $1842 m0 *1 29.375,74.75
X$1842 165 166 167 231 168 232 257 258 cell_2rw
* cell instance $1843 r0 *1 29.375,74.75
X$1843 165 166 167 230 168 229 257 258 cell_2rw
* cell instance $1844 m0 *1 29.375,77.74
X$1844 165 166 167 227 168 228 257 258 cell_2rw
* cell instance $1845 m0 *1 29.375,80.73
X$1845 165 166 167 233 168 236 257 258 cell_2rw
* cell instance $1846 r0 *1 29.375,77.74
X$1846 165 166 167 237 168 238 257 258 cell_2rw
* cell instance $1847 r0 *1 29.375,80.73
X$1847 165 166 167 235 168 234 257 258 cell_2rw
* cell instance $1848 m0 *1 29.375,83.72
X$1848 165 166 167 240 168 242 257 258 cell_2rw
* cell instance $1849 r0 *1 29.375,83.72
X$1849 165 166 167 239 168 241 257 258 cell_2rw
* cell instance $1850 m0 *1 29.375,86.71
X$1850 165 166 167 244 168 243 257 258 cell_2rw
* cell instance $1851 r0 *1 29.375,86.71
X$1851 165 166 167 245 168 247 257 258 cell_2rw
* cell instance $1852 m0 *1 29.375,89.7
X$1852 165 166 167 250 168 249 257 258 cell_2rw
* cell instance $1853 r0 *1 29.375,89.7
X$1853 165 166 167 246 168 248 257 258 cell_2rw
* cell instance $1854 m0 *1 29.375,92.69
X$1854 165 166 167 253 168 256 257 258 cell_2rw
* cell instance $1855 m0 *1 29.375,95.68
X$1855 165 166 167 251 168 252 257 258 cell_2rw
* cell instance $1856 r0 *1 29.375,92.69
X$1856 165 166 167 255 168 254 257 258 cell_2rw
* cell instance $1857 r0 *1 30.55,47.84
X$1857 169 170 171 199 172 201 257 258 cell_2rw
* cell instance $1858 m0 *1 30.55,50.83
X$1858 169 170 171 195 172 197 257 258 cell_2rw
* cell instance $1859 r0 *1 30.55,50.83
X$1859 169 170 171 202 172 194 257 258 cell_2rw
* cell instance $1860 m0 *1 30.55,53.82
X$1860 169 170 171 198 172 193 257 258 cell_2rw
* cell instance $1861 r0 *1 30.55,53.82
X$1861 169 170 171 196 172 200 257 258 cell_2rw
* cell instance $1862 m0 *1 30.55,56.81
X$1862 169 170 171 203 172 207 257 258 cell_2rw
* cell instance $1863 r0 *1 30.55,56.81
X$1863 169 170 171 206 172 208 257 258 cell_2rw
* cell instance $1864 m0 *1 30.55,59.8
X$1864 169 170 171 205 172 204 257 258 cell_2rw
* cell instance $1865 r0 *1 30.55,59.8
X$1865 169 170 171 214 172 213 257 258 cell_2rw
* cell instance $1866 m0 *1 30.55,62.79
X$1866 169 170 171 212 172 211 257 258 cell_2rw
* cell instance $1867 m0 *1 30.55,65.78
X$1867 169 170 171 219 172 217 257 258 cell_2rw
* cell instance $1868 r0 *1 30.55,62.79
X$1868 169 170 171 210 172 209 257 258 cell_2rw
* cell instance $1869 m0 *1 30.55,68.77
X$1869 169 170 171 218 172 220 257 258 cell_2rw
* cell instance $1870 r0 *1 30.55,65.78
X$1870 169 170 171 216 172 215 257 258 cell_2rw
* cell instance $1871 r0 *1 30.55,68.77
X$1871 169 170 171 224 172 223 257 258 cell_2rw
* cell instance $1872 m0 *1 30.55,71.76
X$1872 169 170 171 221 172 222 257 258 cell_2rw
* cell instance $1873 r0 *1 30.55,71.76
X$1873 169 170 171 226 172 225 257 258 cell_2rw
* cell instance $1874 m0 *1 30.55,74.75
X$1874 169 170 171 231 172 232 257 258 cell_2rw
* cell instance $1875 r0 *1 30.55,74.75
X$1875 169 170 171 230 172 229 257 258 cell_2rw
* cell instance $1876 m0 *1 30.55,77.74
X$1876 169 170 171 227 172 228 257 258 cell_2rw
* cell instance $1877 r0 *1 30.55,77.74
X$1877 169 170 171 237 172 238 257 258 cell_2rw
* cell instance $1878 m0 *1 30.55,80.73
X$1878 169 170 171 233 172 236 257 258 cell_2rw
* cell instance $1879 r0 *1 30.55,80.73
X$1879 169 170 171 235 172 234 257 258 cell_2rw
* cell instance $1880 m0 *1 30.55,83.72
X$1880 169 170 171 240 172 242 257 258 cell_2rw
* cell instance $1881 r0 *1 30.55,83.72
X$1881 169 170 171 239 172 241 257 258 cell_2rw
* cell instance $1882 m0 *1 30.55,86.71
X$1882 169 170 171 244 172 243 257 258 cell_2rw
* cell instance $1883 r0 *1 30.55,86.71
X$1883 169 170 171 245 172 247 257 258 cell_2rw
* cell instance $1884 m0 *1 30.55,89.7
X$1884 169 170 171 250 172 249 257 258 cell_2rw
* cell instance $1885 m0 *1 30.55,92.69
X$1885 169 170 171 253 172 256 257 258 cell_2rw
* cell instance $1886 r0 *1 30.55,89.7
X$1886 169 170 171 246 172 248 257 258 cell_2rw
* cell instance $1887 r0 *1 30.55,92.69
X$1887 169 170 171 255 172 254 257 258 cell_2rw
* cell instance $1888 m0 *1 30.55,95.68
X$1888 169 170 171 251 172 252 257 258 cell_2rw
* cell instance $1889 r0 *1 31.725,47.84
X$1889 173 174 175 199 176 201 257 258 cell_2rw
* cell instance $1890 m0 *1 31.725,50.83
X$1890 173 174 175 195 176 197 257 258 cell_2rw
* cell instance $1891 r0 *1 31.725,50.83
X$1891 173 174 175 202 176 194 257 258 cell_2rw
* cell instance $1892 m0 *1 31.725,53.82
X$1892 173 174 175 198 176 193 257 258 cell_2rw
* cell instance $1893 r0 *1 31.725,53.82
X$1893 173 174 175 196 176 200 257 258 cell_2rw
* cell instance $1894 m0 *1 31.725,56.81
X$1894 173 174 175 203 176 207 257 258 cell_2rw
* cell instance $1895 r0 *1 31.725,56.81
X$1895 173 174 175 206 176 208 257 258 cell_2rw
* cell instance $1896 m0 *1 31.725,59.8
X$1896 173 174 175 205 176 204 257 258 cell_2rw
* cell instance $1897 r0 *1 31.725,59.8
X$1897 173 174 175 214 176 213 257 258 cell_2rw
* cell instance $1898 m0 *1 31.725,62.79
X$1898 173 174 175 212 176 211 257 258 cell_2rw
* cell instance $1899 r0 *1 31.725,62.79
X$1899 173 174 175 210 176 209 257 258 cell_2rw
* cell instance $1900 m0 *1 31.725,65.78
X$1900 173 174 175 219 176 217 257 258 cell_2rw
* cell instance $1901 r0 *1 31.725,65.78
X$1901 173 174 175 216 176 215 257 258 cell_2rw
* cell instance $1902 m0 *1 31.725,68.77
X$1902 173 174 175 218 176 220 257 258 cell_2rw
* cell instance $1903 m0 *1 31.725,71.76
X$1903 173 174 175 221 176 222 257 258 cell_2rw
* cell instance $1904 r0 *1 31.725,68.77
X$1904 173 174 175 224 176 223 257 258 cell_2rw
* cell instance $1905 m0 *1 31.725,74.75
X$1905 173 174 175 231 176 232 257 258 cell_2rw
* cell instance $1906 r0 *1 31.725,71.76
X$1906 173 174 175 226 176 225 257 258 cell_2rw
* cell instance $1907 r0 *1 31.725,74.75
X$1907 173 174 175 230 176 229 257 258 cell_2rw
* cell instance $1908 m0 *1 31.725,77.74
X$1908 173 174 175 227 176 228 257 258 cell_2rw
* cell instance $1909 r0 *1 31.725,77.74
X$1909 173 174 175 237 176 238 257 258 cell_2rw
* cell instance $1910 m0 *1 31.725,80.73
X$1910 173 174 175 233 176 236 257 258 cell_2rw
* cell instance $1911 r0 *1 31.725,80.73
X$1911 173 174 175 235 176 234 257 258 cell_2rw
* cell instance $1912 m0 *1 31.725,83.72
X$1912 173 174 175 240 176 242 257 258 cell_2rw
* cell instance $1913 r0 *1 31.725,83.72
X$1913 173 174 175 239 176 241 257 258 cell_2rw
* cell instance $1914 m0 *1 31.725,86.71
X$1914 173 174 175 244 176 243 257 258 cell_2rw
* cell instance $1915 r0 *1 31.725,86.71
X$1915 173 174 175 245 176 247 257 258 cell_2rw
* cell instance $1916 m0 *1 31.725,89.7
X$1916 173 174 175 250 176 249 257 258 cell_2rw
* cell instance $1917 r0 *1 31.725,89.7
X$1917 173 174 175 246 176 248 257 258 cell_2rw
* cell instance $1918 m0 *1 31.725,92.69
X$1918 173 174 175 253 176 256 257 258 cell_2rw
* cell instance $1919 r0 *1 31.725,92.69
X$1919 173 174 175 255 176 254 257 258 cell_2rw
* cell instance $1920 m0 *1 31.725,95.68
X$1920 173 174 175 251 176 252 257 258 cell_2rw
* cell instance $1921 r0 *1 32.9,47.84
X$1921 177 178 179 199 180 201 257 258 cell_2rw
* cell instance $1922 m0 *1 32.9,50.83
X$1922 177 178 179 195 180 197 257 258 cell_2rw
* cell instance $1923 r0 *1 32.9,50.83
X$1923 177 178 179 202 180 194 257 258 cell_2rw
* cell instance $1924 m0 *1 32.9,53.82
X$1924 177 178 179 198 180 193 257 258 cell_2rw
* cell instance $1925 r0 *1 32.9,53.82
X$1925 177 178 179 196 180 200 257 258 cell_2rw
* cell instance $1926 m0 *1 32.9,56.81
X$1926 177 178 179 203 180 207 257 258 cell_2rw
* cell instance $1927 r0 *1 32.9,56.81
X$1927 177 178 179 206 180 208 257 258 cell_2rw
* cell instance $1928 m0 *1 32.9,59.8
X$1928 177 178 179 205 180 204 257 258 cell_2rw
* cell instance $1929 r0 *1 32.9,59.8
X$1929 177 178 179 214 180 213 257 258 cell_2rw
* cell instance $1930 m0 *1 32.9,62.79
X$1930 177 178 179 212 180 211 257 258 cell_2rw
* cell instance $1931 r0 *1 32.9,62.79
X$1931 177 178 179 210 180 209 257 258 cell_2rw
* cell instance $1932 m0 *1 32.9,65.78
X$1932 177 178 179 219 180 217 257 258 cell_2rw
* cell instance $1933 r0 *1 32.9,65.78
X$1933 177 178 179 216 180 215 257 258 cell_2rw
* cell instance $1934 m0 *1 32.9,68.77
X$1934 177 178 179 218 180 220 257 258 cell_2rw
* cell instance $1935 m0 *1 32.9,71.76
X$1935 177 178 179 221 180 222 257 258 cell_2rw
* cell instance $1936 r0 *1 32.9,68.77
X$1936 177 178 179 224 180 223 257 258 cell_2rw
* cell instance $1937 m0 *1 32.9,74.75
X$1937 177 178 179 231 180 232 257 258 cell_2rw
* cell instance $1938 r0 *1 32.9,71.76
X$1938 177 178 179 226 180 225 257 258 cell_2rw
* cell instance $1939 r0 *1 32.9,74.75
X$1939 177 178 179 230 180 229 257 258 cell_2rw
* cell instance $1940 m0 *1 32.9,77.74
X$1940 177 178 179 227 180 228 257 258 cell_2rw
* cell instance $1941 r0 *1 32.9,77.74
X$1941 177 178 179 237 180 238 257 258 cell_2rw
* cell instance $1942 m0 *1 32.9,80.73
X$1942 177 178 179 233 180 236 257 258 cell_2rw
* cell instance $1943 r0 *1 32.9,80.73
X$1943 177 178 179 235 180 234 257 258 cell_2rw
* cell instance $1944 m0 *1 32.9,83.72
X$1944 177 178 179 240 180 242 257 258 cell_2rw
* cell instance $1945 r0 *1 32.9,83.72
X$1945 177 178 179 239 180 241 257 258 cell_2rw
* cell instance $1946 m0 *1 32.9,86.71
X$1946 177 178 179 244 180 243 257 258 cell_2rw
* cell instance $1947 m0 *1 32.9,89.7
X$1947 177 178 179 250 180 249 257 258 cell_2rw
* cell instance $1948 r0 *1 32.9,86.71
X$1948 177 178 179 245 180 247 257 258 cell_2rw
* cell instance $1949 r0 *1 32.9,89.7
X$1949 177 178 179 246 180 248 257 258 cell_2rw
* cell instance $1950 m0 *1 32.9,92.69
X$1950 177 178 179 253 180 256 257 258 cell_2rw
* cell instance $1951 r0 *1 32.9,92.69
X$1951 177 178 179 255 180 254 257 258 cell_2rw
* cell instance $1952 m0 *1 32.9,95.68
X$1952 177 178 179 251 180 252 257 258 cell_2rw
* cell instance $1953 r0 *1 34.075,47.84
X$1953 181 182 183 199 184 201 257 258 cell_2rw
* cell instance $1954 m0 *1 34.075,50.83
X$1954 181 182 183 195 184 197 257 258 cell_2rw
* cell instance $1955 r0 *1 34.075,50.83
X$1955 181 182 183 202 184 194 257 258 cell_2rw
* cell instance $1956 m0 *1 34.075,53.82
X$1956 181 182 183 198 184 193 257 258 cell_2rw
* cell instance $1957 r0 *1 34.075,53.82
X$1957 181 182 183 196 184 200 257 258 cell_2rw
* cell instance $1958 m0 *1 34.075,56.81
X$1958 181 182 183 203 184 207 257 258 cell_2rw
* cell instance $1959 r0 *1 34.075,56.81
X$1959 181 182 183 206 184 208 257 258 cell_2rw
* cell instance $1960 m0 *1 34.075,59.8
X$1960 181 182 183 205 184 204 257 258 cell_2rw
* cell instance $1961 m0 *1 34.075,62.79
X$1961 181 182 183 212 184 211 257 258 cell_2rw
* cell instance $1962 r0 *1 34.075,59.8
X$1962 181 182 183 214 184 213 257 258 cell_2rw
* cell instance $1963 r0 *1 34.075,62.79
X$1963 181 182 183 210 184 209 257 258 cell_2rw
* cell instance $1964 m0 *1 34.075,65.78
X$1964 181 182 183 219 184 217 257 258 cell_2rw
* cell instance $1965 r0 *1 34.075,65.78
X$1965 181 182 183 216 184 215 257 258 cell_2rw
* cell instance $1966 m0 *1 34.075,68.77
X$1966 181 182 183 218 184 220 257 258 cell_2rw
* cell instance $1967 r0 *1 34.075,68.77
X$1967 181 182 183 224 184 223 257 258 cell_2rw
* cell instance $1968 m0 *1 34.075,71.76
X$1968 181 182 183 221 184 222 257 258 cell_2rw
* cell instance $1969 r0 *1 34.075,71.76
X$1969 181 182 183 226 184 225 257 258 cell_2rw
* cell instance $1970 m0 *1 34.075,74.75
X$1970 181 182 183 231 184 232 257 258 cell_2rw
* cell instance $1971 r0 *1 34.075,74.75
X$1971 181 182 183 230 184 229 257 258 cell_2rw
* cell instance $1972 m0 *1 34.075,77.74
X$1972 181 182 183 227 184 228 257 258 cell_2rw
* cell instance $1973 r0 *1 34.075,77.74
X$1973 181 182 183 237 184 238 257 258 cell_2rw
* cell instance $1974 m0 *1 34.075,80.73
X$1974 181 182 183 233 184 236 257 258 cell_2rw
* cell instance $1975 r0 *1 34.075,80.73
X$1975 181 182 183 235 184 234 257 258 cell_2rw
* cell instance $1976 m0 *1 34.075,83.72
X$1976 181 182 183 240 184 242 257 258 cell_2rw
* cell instance $1977 r0 *1 34.075,83.72
X$1977 181 182 183 239 184 241 257 258 cell_2rw
* cell instance $1978 m0 *1 34.075,86.71
X$1978 181 182 183 244 184 243 257 258 cell_2rw
* cell instance $1979 m0 *1 34.075,89.7
X$1979 181 182 183 250 184 249 257 258 cell_2rw
* cell instance $1980 r0 *1 34.075,86.71
X$1980 181 182 183 245 184 247 257 258 cell_2rw
* cell instance $1981 r0 *1 34.075,89.7
X$1981 181 182 183 246 184 248 257 258 cell_2rw
* cell instance $1982 m0 *1 34.075,92.69
X$1982 181 182 183 253 184 256 257 258 cell_2rw
* cell instance $1983 r0 *1 34.075,92.69
X$1983 181 182 183 255 184 254 257 258 cell_2rw
* cell instance $1984 m0 *1 34.075,95.68
X$1984 181 182 183 251 184 252 257 258 cell_2rw
* cell instance $1985 r0 *1 35.25,47.84
X$1985 185 186 187 199 188 201 257 258 cell_2rw
* cell instance $1986 m0 *1 35.25,50.83
X$1986 185 186 187 195 188 197 257 258 cell_2rw
* cell instance $1987 r0 *1 35.25,50.83
X$1987 185 186 187 202 188 194 257 258 cell_2rw
* cell instance $1988 m0 *1 35.25,53.82
X$1988 185 186 187 198 188 193 257 258 cell_2rw
* cell instance $1989 m0 *1 35.25,56.81
X$1989 185 186 187 203 188 207 257 258 cell_2rw
* cell instance $1990 r0 *1 35.25,53.82
X$1990 185 186 187 196 188 200 257 258 cell_2rw
* cell instance $1991 r0 *1 35.25,56.81
X$1991 185 186 187 206 188 208 257 258 cell_2rw
* cell instance $1992 m0 *1 35.25,59.8
X$1992 185 186 187 205 188 204 257 258 cell_2rw
* cell instance $1993 r0 *1 35.25,59.8
X$1993 185 186 187 214 188 213 257 258 cell_2rw
* cell instance $1994 m0 *1 35.25,62.79
X$1994 185 186 187 212 188 211 257 258 cell_2rw
* cell instance $1995 r0 *1 35.25,62.79
X$1995 185 186 187 210 188 209 257 258 cell_2rw
* cell instance $1996 m0 *1 35.25,65.78
X$1996 185 186 187 219 188 217 257 258 cell_2rw
* cell instance $1997 r0 *1 35.25,65.78
X$1997 185 186 187 216 188 215 257 258 cell_2rw
* cell instance $1998 m0 *1 35.25,68.77
X$1998 185 186 187 218 188 220 257 258 cell_2rw
* cell instance $1999 m0 *1 35.25,71.76
X$1999 185 186 187 221 188 222 257 258 cell_2rw
* cell instance $2000 r0 *1 35.25,68.77
X$2000 185 186 187 224 188 223 257 258 cell_2rw
* cell instance $2001 r0 *1 35.25,71.76
X$2001 185 186 187 226 188 225 257 258 cell_2rw
* cell instance $2002 m0 *1 35.25,74.75
X$2002 185 186 187 231 188 232 257 258 cell_2rw
* cell instance $2003 m0 *1 35.25,77.74
X$2003 185 186 187 227 188 228 257 258 cell_2rw
* cell instance $2004 r0 *1 35.25,74.75
X$2004 185 186 187 230 188 229 257 258 cell_2rw
* cell instance $2005 r0 *1 35.25,77.74
X$2005 185 186 187 237 188 238 257 258 cell_2rw
* cell instance $2006 m0 *1 35.25,80.73
X$2006 185 186 187 233 188 236 257 258 cell_2rw
* cell instance $2007 r0 *1 35.25,80.73
X$2007 185 186 187 235 188 234 257 258 cell_2rw
* cell instance $2008 m0 *1 35.25,83.72
X$2008 185 186 187 240 188 242 257 258 cell_2rw
* cell instance $2009 r0 *1 35.25,83.72
X$2009 185 186 187 239 188 241 257 258 cell_2rw
* cell instance $2010 m0 *1 35.25,86.71
X$2010 185 186 187 244 188 243 257 258 cell_2rw
* cell instance $2011 r0 *1 35.25,86.71
X$2011 185 186 187 245 188 247 257 258 cell_2rw
* cell instance $2012 m0 *1 35.25,89.7
X$2012 185 186 187 250 188 249 257 258 cell_2rw
* cell instance $2013 r0 *1 35.25,89.7
X$2013 185 186 187 246 188 248 257 258 cell_2rw
* cell instance $2014 m0 *1 35.25,92.69
X$2014 185 186 187 253 188 256 257 258 cell_2rw
* cell instance $2015 m0 *1 35.25,95.68
X$2015 185 186 187 251 188 252 257 258 cell_2rw
* cell instance $2016 r0 *1 35.25,92.69
X$2016 185 186 187 255 188 254 257 258 cell_2rw
* cell instance $2017 r0 *1 36.425,47.84
X$2017 189 190 191 199 192 201 257 258 cell_2rw
* cell instance $2018 m0 *1 36.425,50.83
X$2018 189 190 191 195 192 197 257 258 cell_2rw
* cell instance $2019 r0 *1 36.425,50.83
X$2019 189 190 191 202 192 194 257 258 cell_2rw
* cell instance $2020 m0 *1 36.425,53.82
X$2020 189 190 191 198 192 193 257 258 cell_2rw
* cell instance $2021 r0 *1 36.425,53.82
X$2021 189 190 191 196 192 200 257 258 cell_2rw
* cell instance $2022 m0 *1 36.425,56.81
X$2022 189 190 191 203 192 207 257 258 cell_2rw
* cell instance $2023 m0 *1 36.425,59.8
X$2023 189 190 191 205 192 204 257 258 cell_2rw
* cell instance $2024 r0 *1 36.425,56.81
X$2024 189 190 191 206 192 208 257 258 cell_2rw
* cell instance $2025 r0 *1 36.425,59.8
X$2025 189 190 191 214 192 213 257 258 cell_2rw
* cell instance $2026 m0 *1 36.425,62.79
X$2026 189 190 191 212 192 211 257 258 cell_2rw
* cell instance $2027 r0 *1 36.425,62.79
X$2027 189 190 191 210 192 209 257 258 cell_2rw
* cell instance $2028 m0 *1 36.425,65.78
X$2028 189 190 191 219 192 217 257 258 cell_2rw
* cell instance $2029 m0 *1 36.425,68.77
X$2029 189 190 191 218 192 220 257 258 cell_2rw
* cell instance $2030 r0 *1 36.425,65.78
X$2030 189 190 191 216 192 215 257 258 cell_2rw
* cell instance $2031 r0 *1 36.425,68.77
X$2031 189 190 191 224 192 223 257 258 cell_2rw
* cell instance $2032 m0 *1 36.425,71.76
X$2032 189 190 191 221 192 222 257 258 cell_2rw
* cell instance $2033 r0 *1 36.425,71.76
X$2033 189 190 191 226 192 225 257 258 cell_2rw
* cell instance $2034 m0 *1 36.425,74.75
X$2034 189 190 191 231 192 232 257 258 cell_2rw
* cell instance $2035 r0 *1 36.425,74.75
X$2035 189 190 191 230 192 229 257 258 cell_2rw
* cell instance $2036 m0 *1 36.425,77.74
X$2036 189 190 191 227 192 228 257 258 cell_2rw
* cell instance $2037 r0 *1 36.425,77.74
X$2037 189 190 191 237 192 238 257 258 cell_2rw
* cell instance $2038 m0 *1 36.425,80.73
X$2038 189 190 191 233 192 236 257 258 cell_2rw
* cell instance $2039 r0 *1 36.425,80.73
X$2039 189 190 191 235 192 234 257 258 cell_2rw
* cell instance $2040 m0 *1 36.425,83.72
X$2040 189 190 191 240 192 242 257 258 cell_2rw
* cell instance $2041 r0 *1 36.425,83.72
X$2041 189 190 191 239 192 241 257 258 cell_2rw
* cell instance $2042 m0 *1 36.425,86.71
X$2042 189 190 191 244 192 243 257 258 cell_2rw
* cell instance $2043 r0 *1 36.425,86.71
X$2043 189 190 191 245 192 247 257 258 cell_2rw
* cell instance $2044 m0 *1 36.425,89.7
X$2044 189 190 191 250 192 249 257 258 cell_2rw
* cell instance $2045 r0 *1 36.425,89.7
X$2045 189 190 191 246 192 248 257 258 cell_2rw
* cell instance $2046 m0 *1 36.425,92.69
X$2046 189 190 191 253 192 256 257 258 cell_2rw
* cell instance $2047 r0 *1 36.425,92.69
X$2047 189 190 191 255 192 254 257 258 cell_2rw
* cell instance $2048 m0 *1 36.425,95.68
X$2048 189 190 191 251 192 252 257 258 cell_2rw
.ENDS custom_sram_1r1w_32_256_freepdk45_bitcell_array

* cell dummy_cell_2rw
* pin wl1
* pin wl0
* pin vdd
* pin gnd
.SUBCKT dummy_cell_2rw 1 9 11 12
* net 1 wl1
* net 9 wl0
* net 11 vdd
* net 12 gnd
* device instance $1 r0 *1 0.4925,1.2075 PMOS_VTG
M$1 10 3 11 11 PMOS_VTG L=0.05U W=0.09U AS=0.00945P AD=0.0063P PS=0.39U PD=0.23U
* device instance $2 r0 *1 0.6825,1.2075 PMOS_VTG
M$2 11 10 3 11 PMOS_VTG L=0.05U W=0.09U AS=0.0063P AD=0.00945P PS=0.23U PD=0.39U
* device instance $3 r0 *1 0.2875,0.69 NMOS_VTG
M$3 10 9 7 12 NMOS_VTG L=0.05U W=0.135U AS=0.0141375P AD=0.014175P PS=0.36U
+ PD=0.48U
* device instance $4 r0 *1 0.4925,0.655 NMOS_VTG
M$4 10 3 12 12 NMOS_VTG L=0.05U W=0.205U AS=0.0141375P AD=0.01435P PS=0.36U
+ PD=0.345U
* device instance $5 r0 *1 0.6825,0.655 NMOS_VTG
M$5 12 10 3 12 NMOS_VTG L=0.05U W=0.205U AS=0.01435P AD=0.0141375P PS=0.345U
+ PD=0.36U
* device instance $6 r0 *1 0.8875,0.69 NMOS_VTG
M$6 3 9 8 12 NMOS_VTG L=0.05U W=0.135U AS=0.0141375P AD=0.014175P PS=0.36U
+ PD=0.48U
* device instance $7 r0 *1 0.3025,0.3225 NMOS_VTG
M$7 2 1 5 12 NMOS_VTG L=0.05U W=0.18U AS=0.02025P AD=0.0126P PS=0.585U PD=0.32U
* device instance $8 r0 *1 0.4925,0.3225 NMOS_VTG
M$8 5 3 12 12 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.0126P PS=0.32U PD=0.32U
* device instance $9 r0 *1 0.6825,0.3225 NMOS_VTG
M$9 12 10 6 12 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.0126P PS=0.32U PD=0.32U
* device instance $10 r0 *1 0.8725,0.3225 NMOS_VTG
M$10 6 1 4 12 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.02025P PS=0.32U PD=0.585U
.ENDS dummy_cell_2rw

* cell replica_cell_2rw
* pin bl0
* pin bl1
* pin br1
* pin wl1
* pin br0
* pin wl0
* pin vdd
* pin gnd
.SUBCKT replica_cell_2rw 1 2 3 4 7 8 10 11
* net 1 bl0
* net 2 bl1
* net 3 br1
* net 4 wl1
* net 7 br0
* net 8 wl0
* net 10 vdd
* net 11 gnd
* device instance $1 r0 *1 0.4925,1.2075 PMOS_VTG
M$1 9 10 10 10 PMOS_VTG L=0.05U W=0.09U AS=0.00945P AD=0.0063P PS=0.39U PD=0.23U
* device instance $2 r0 *1 0.6825,1.2075 PMOS_VTG
M$2 10 9 10 10 PMOS_VTG L=0.05U W=0.09U AS=0.0063P AD=0.00945P PS=0.23U PD=0.39U
* device instance $3 r0 *1 0.2875,0.69 NMOS_VTG
M$3 9 8 1 11 NMOS_VTG L=0.05U W=0.135U AS=0.0141375P AD=0.014175P PS=0.36U
+ PD=0.48U
* device instance $4 r0 *1 0.4925,0.655 NMOS_VTG
M$4 9 10 11 11 NMOS_VTG L=0.05U W=0.205U AS=0.0141375P AD=0.01435P PS=0.36U
+ PD=0.345U
* device instance $5 r0 *1 0.6825,0.655 NMOS_VTG
M$5 11 9 10 11 NMOS_VTG L=0.05U W=0.205U AS=0.01435P AD=0.0141375P PS=0.345U
+ PD=0.36U
* device instance $6 r0 *1 0.8875,0.69 NMOS_VTG
M$6 10 8 7 11 NMOS_VTG L=0.05U W=0.135U AS=0.0141375P AD=0.014175P PS=0.36U
+ PD=0.48U
* device instance $7 r0 *1 0.3025,0.3225 NMOS_VTG
M$7 2 4 5 11 NMOS_VTG L=0.05U W=0.18U AS=0.02025P AD=0.0126P PS=0.585U PD=0.32U
* device instance $8 r0 *1 0.4925,0.3225 NMOS_VTG
M$8 5 10 11 11 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.0126P PS=0.32U PD=0.32U
* device instance $9 r0 *1 0.6825,0.3225 NMOS_VTG
M$9 11 9 6 11 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.0126P PS=0.32U PD=0.32U
* device instance $10 r0 *1 0.8725,0.3225 NMOS_VTG
M$10 6 4 3 11 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.02025P PS=0.32U PD=0.585U
.ENDS replica_cell_2rw

* cell cell_2rw
* pin bl0
* pin bl1
* pin br1
* pin wl1
* pin br0
* pin wl0
* pin vdd
* pin gnd
.SUBCKT cell_2rw 1 2 3 4 8 9 11 12
* net 1 bl0
* net 2 bl1
* net 3 br1
* net 4 wl1
* net 8 br0
* net 9 wl0
* net 11 vdd
* net 12 gnd
* device instance $1 r0 *1 0.4925,1.2075 PMOS_VTG
M$1 10 5 11 11 PMOS_VTG L=0.05U W=0.09U AS=0.00945P AD=0.0063P PS=0.39U PD=0.23U
* device instance $2 r0 *1 0.6825,1.2075 PMOS_VTG
M$2 11 10 5 11 PMOS_VTG L=0.05U W=0.09U AS=0.0063P AD=0.00945P PS=0.23U PD=0.39U
* device instance $3 r0 *1 0.2875,0.69 NMOS_VTG
M$3 10 9 1 12 NMOS_VTG L=0.05U W=0.135U AS=0.0141375P AD=0.014175P PS=0.36U
+ PD=0.48U
* device instance $4 r0 *1 0.4925,0.655 NMOS_VTG
M$4 10 5 12 12 NMOS_VTG L=0.05U W=0.205U AS=0.0141375P AD=0.01435P PS=0.36U
+ PD=0.345U
* device instance $5 r0 *1 0.6825,0.655 NMOS_VTG
M$5 12 10 5 12 NMOS_VTG L=0.05U W=0.205U AS=0.01435P AD=0.0141375P PS=0.345U
+ PD=0.36U
* device instance $6 r0 *1 0.8875,0.69 NMOS_VTG
M$6 5 9 8 12 NMOS_VTG L=0.05U W=0.135U AS=0.0141375P AD=0.014175P PS=0.36U
+ PD=0.48U
* device instance $7 r0 *1 0.3025,0.3225 NMOS_VTG
M$7 2 4 6 12 NMOS_VTG L=0.05U W=0.18U AS=0.02025P AD=0.0126P PS=0.585U PD=0.32U
* device instance $8 r0 *1 0.4925,0.3225 NMOS_VTG
M$8 6 5 12 12 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.0126P PS=0.32U PD=0.32U
* device instance $9 r0 *1 0.6825,0.3225 NMOS_VTG
M$9 12 10 7 12 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.0126P PS=0.32U PD=0.32U
* device instance $10 r0 *1 0.8725,0.3225 NMOS_VTG
M$10 7 4 3 12 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.02025P PS=0.32U PD=0.585U
.ENDS cell_2rw
